-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 22.03.2012 9:17:45
-- Module Name : usrif_cfg
--
-- Description : ����� ���������� ����������
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package usrif_cfg is

constant C_HSCAM_USRIF : string:="FTDI";

end usrif_cfg;

