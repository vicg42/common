-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 25.11.2008 18:38
-- Module Name : vsobel_main_tb
--
-- ����������/�������� :
--    �������� ������
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_textio.all;

use work.vicg_common_pkg.all;

library std;
use std.textio.all;

library unisim;
use unisim.vcomponents.all;

entity vsobel_main_tb is
end vsobel_main_tb;

architecture behavior of vsobel_main_tb is

constant i_clk_period : TIME := 6.6 ns; --150MHz

----//�������� �������� - tst.png
--type TImageTst  is array (0 to (8*17)-1) of std_logic_vector (31 downto 0);
--constant C_TST_IMAGE : TImageTst:=(
----//Y0
--(CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#178#, 8)&CONV_STD_LOGIC_VECTOR(10#163#, 8)&CONV_STD_LOGIC_VECTOR(10#096#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#117#, 8)&CONV_STD_LOGIC_VECTOR(10#157#, 8)&CONV_STD_LOGIC_VECTOR(10#160#, 8)&CONV_STD_LOGIC_VECTOR(10#161#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y1
--(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#053#, 8)&CONV_STD_LOGIC_VECTOR(10#086#, 8)&CONV_STD_LOGIC_VECTOR(10#047#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#036#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#172#, 8)&CONV_STD_LOGIC_VECTOR(10#174#, 8)&CONV_STD_LOGIC_VECTOR(10#119#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#107#, 8)&CONV_STD_LOGIC_VECTOR(10#152#, 8)&CONV_STD_LOGIC_VECTOR(10#157#, 8)&CONV_STD_LOGIC_VECTOR(10#155#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y2
--(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#135#, 8)&CONV_STD_LOGIC_VECTOR(10#077#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#179#, 8)&CONV_STD_LOGIC_VECTOR(10#234#, 8)&CONV_STD_LOGIC_VECTOR(10#190#, 8)&CONV_STD_LOGIC_VECTOR(10#152#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#068#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#179#, 8)&CONV_STD_LOGIC_VECTOR(10#195#, 8)&CONV_STD_LOGIC_VECTOR(10#159#, 8)&CONV_STD_LOGIC_VECTOR(10#045#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#076#, 8)&CONV_STD_LOGIC_VECTOR(10#132#, 8)&CONV_STD_LOGIC_VECTOR(10#154#, 8)&CONV_STD_LOGIC_VECTOR(10#161#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y3
--(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#227#, 8)&CONV_STD_LOGIC_VECTOR(10#107#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#032#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#242#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#243#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#009#, 8)&CONV_STD_LOGIC_VECTOR(10#007#, 8)&CONV_STD_LOGIC_VECTOR(10#063#, 8)&CONV_STD_LOGIC_VECTOR(10#169#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#219#, 8)&CONV_STD_LOGIC_VECTOR(10#235#, 8)&CONV_STD_LOGIC_VECTOR(10#211#, 8)&CONV_STD_LOGIC_VECTOR(10#087#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#064#, 8)&CONV_STD_LOGIC_VECTOR(10#136#, 8)&CONV_STD_LOGIC_VECTOR(10#187#, 8)&CONV_STD_LOGIC_VECTOR(10#207#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y4
--(CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#191#, 8)&CONV_STD_LOGIC_VECTOR(10#074#, 8)&CONV_STD_LOGIC_VECTOR(10#049#, 8)&CONV_STD_LOGIC_VECTOR(10#058#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#247#, 8)&CONV_STD_LOGIC_VECTOR(10#230#, 8)&CONV_STD_LOGIC_VECTOR(10#248#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#053#, 8)&CONV_STD_LOGIC_VECTOR(10#164#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#247#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)&CONV_STD_LOGIC_VECTOR(10#119#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#067#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y5
--(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#097#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#043#, 8)&CONV_STD_LOGIC_VECTOR(10#053#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#243#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#217#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#074#, 8)&CONV_STD_LOGIC_VECTOR(10#143#, 8)&CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#245#, 8)&CONV_STD_LOGIC_VECTOR(10#248#, 8)&CONV_STD_LOGIC_VECTOR(10#245#, 8)&CONV_STD_LOGIC_VECTOR(10#148#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#058#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#244#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y6
--(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#047#, 8)&CONV_STD_LOGIC_VECTOR(10#042#, 8)&CONV_STD_LOGIC_VECTOR(10#077#, 8)&CONV_STD_LOGIC_VECTOR(10#055#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#238#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)&CONV_STD_LOGIC_VECTOR(10#157#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#162#, 8)&CONV_STD_LOGIC_VECTOR(10#214#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#249#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)&CONV_STD_LOGIC_VECTOR(10#253#, 8)&CONV_STD_LOGIC_VECTOR(10#200#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#050#, 8)&CONV_STD_LOGIC_VECTOR(10#139#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#253#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y7
--(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#065#, 8)&CONV_STD_LOGIC_VECTOR(10#127#, 8)&CONV_STD_LOGIC_VECTOR(10#172#, 8)&CONV_STD_LOGIC_VECTOR(10#106#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#249#, 8)&CONV_STD_LOGIC_VECTOR(10#251#, 8)&CONV_STD_LOGIC_VECTOR(10#205#, 8)&CONV_STD_LOGIC_VECTOR(10#091#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#221#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)&CONV_STD_LOGIC_VECTOR(10#247#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#239#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#048#, 8)&CONV_STD_LOGIC_VECTOR(10#120#, 8)&CONV_STD_LOGIC_VECTOR(10#216#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y8
--(CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#009#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#159#, 8)&CONV_STD_LOGIC_VECTOR(10#199#, 8)&CONV_STD_LOGIC_VECTOR(10#198#, 8)&CONV_STD_LOGIC_VECTOR(10#107#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#226#, 8)&CONV_STD_LOGIC_VECTOR(10#143#, 8)&CONV_STD_LOGIC_VECTOR(10#105#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#228#, 8)&CONV_STD_LOGIC_VECTOR(10#237#, 8)&CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#247#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#239#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)&CONV_STD_LOGIC_VECTOR(10#248#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#125#, 8)&CONV_STD_LOGIC_VECTOR(10#144#, 8)&CONV_STD_LOGIC_VECTOR(10#237#, 8)&CONV_STD_LOGIC_VECTOR(10#252#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y9
--(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#032#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#175#, 8)&CONV_STD_LOGIC_VECTOR(10#165#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#091#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#219#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#127#, 8)&CONV_STD_LOGIC_VECTOR(10#154#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#220#, 8)&CONV_STD_LOGIC_VECTOR(10#235#, 8)&CONV_STD_LOGIC_VECTOR(10#254#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#252#, 8)&CONV_STD_LOGIC_VECTOR(10#253#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#145#, 8)&CONV_STD_LOGIC_VECTOR(10#121#, 8)&CONV_STD_LOGIC_VECTOR(10#211#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y10
--(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#034#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#181#, 8)&CONV_STD_LOGIC_VECTOR(10#184#, 8)&CONV_STD_LOGIC_VECTOR(10#187#, 8)&CONV_STD_LOGIC_VECTOR(10#100#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#183#, 8)&CONV_STD_LOGIC_VECTOR(10#136#, 8)&CONV_STD_LOGIC_VECTOR(10#144#, 8)&CONV_STD_LOGIC_VECTOR(10#183#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#212#, 8)&CONV_STD_LOGIC_VECTOR(10#233#, 8)&CONV_STD_LOGIC_VECTOR(10#249#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#254#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#102#, 8)&CONV_STD_LOGIC_VECTOR(10#084#, 8)&CONV_STD_LOGIC_VECTOR(10#175#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y11
--(CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#038#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#195#, 8)&CONV_STD_LOGIC_VECTOR(10#228#, 8)&CONV_STD_LOGIC_VECTOR(10#218#, 8)&CONV_STD_LOGIC_VECTOR(10#090#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#202#, 8)&CONV_STD_LOGIC_VECTOR(10#204#, 8)&CONV_STD_LOGIC_VECTOR(10#217#, 8)&CONV_STD_LOGIC_VECTOR(10#215#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#220#, 8)&CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#218#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#217#, 8)&CONV_STD_LOGIC_VECTOR(10#216#, 8)&CONV_STD_LOGIC_VECTOR(10#207#, 8)&CONV_STD_LOGIC_VECTOR(10#226#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#131#, 8)&CONV_STD_LOGIC_VECTOR(10#131#, 8)&CONV_STD_LOGIC_VECTOR(10#168#, 8)&CONV_STD_LOGIC_VECTOR(10#198#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y12
--(CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#040#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#140#, 8)&CONV_STD_LOGIC_VECTOR(10#152#, 8)&CONV_STD_LOGIC_VECTOR(10#130#, 8)&CONV_STD_LOGIC_VECTOR(10#039#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#185#, 8)&CONV_STD_LOGIC_VECTOR(10#183#, 8)&CONV_STD_LOGIC_VECTOR(10#174#, 8)&CONV_STD_LOGIC_VECTOR(10#148#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#202#, 8)&CONV_STD_LOGIC_VECTOR(10#206#, 8)&CONV_STD_LOGIC_VECTOR(10#192#, 8)&CONV_STD_LOGIC_VECTOR(10#182#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#172#, 8)&CONV_STD_LOGIC_VECTOR(10#165#, 8)&CONV_STD_LOGIC_VECTOR(10#150#, 8)&CONV_STD_LOGIC_VECTOR(10#175#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#206#, 8)&CONV_STD_LOGIC_VECTOR(10#206#, 8)&CONV_STD_LOGIC_VECTOR(10#187#, 8)&CONV_STD_LOGIC_VECTOR(10#167#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y13
--(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#034#, 8)&CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#046#, 8)&CONV_STD_LOGIC_VECTOR(10#036#, 8)&CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#088#, 8)&CONV_STD_LOGIC_VECTOR(10#067#, 8)&CONV_STD_LOGIC_VECTOR(10#055#, 8)&CONV_STD_LOGIC_VECTOR(10#041#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#146#, 8)&CONV_STD_LOGIC_VECTOR(10#128#, 8)&CONV_STD_LOGIC_VECTOR(10#108#, 8)&CONV_STD_LOGIC_VECTOR(10#094#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#144#, 8)&CONV_STD_LOGIC_VECTOR(10#156#, 8)&CONV_STD_LOGIC_VECTOR(10#143#, 8)&CONV_STD_LOGIC_VECTOR(10#135#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#216#, 8)&CONV_STD_LOGIC_VECTOR(10#224#, 8)&CONV_STD_LOGIC_VECTOR(10#193#, 8)&CONV_STD_LOGIC_VECTOR(10#153#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y14
--(CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#091#, 8)&CONV_STD_LOGIC_VECTOR(10#050#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#128#, 8)&CONV_STD_LOGIC_VECTOR(10#180#, 8)&CONV_STD_LOGIC_VECTOR(10#179#, 8)&CONV_STD_LOGIC_VECTOR(10#151#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#157#, 8)&CONV_STD_LOGIC_VECTOR(10#166#, 8)&CONV_STD_LOGIC_VECTOR(10#129#, 8)&CONV_STD_LOGIC_VECTOR(10#104#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31
--
----//Y15
--(CONV_STD_LOGIC_VECTOR(10#029#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#005#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#041#, 8)&CONV_STD_LOGIC_VECTOR(10#039#, 8)&CONV_STD_LOGIC_VECTOR(10#038#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#075#, 8)&CONV_STD_LOGIC_VECTOR(10#047#, 8)&CONV_STD_LOGIC_VECTOR(10#040#, 8)&CONV_STD_LOGIC_VECTOR(10#041#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#113#, 8)&CONV_STD_LOGIC_VECTOR(10#064#, 8)&CONV_STD_LOGIC_VECTOR(10#071#, 8)&CONV_STD_LOGIC_VECTOR(10#084#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#189#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)&CONV_STD_LOGIC_VECTOR(10#206#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#105#, 8)&CONV_STD_LOGIC_VECTOR(10#114#, 8)&CONV_STD_LOGIC_VECTOR(10#082#, 8)&CONV_STD_LOGIC_VECTOR(10#104#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)),  --//28..31
--
--
----//Y16
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//0..3
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//4..7
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//8..11
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//12..15
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//16..19
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//20..23
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
--(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8))  --//28..31
--
--);

--//�������� �������� - 01g.png (���������� ��� MatLab - 900:915, 900:923)
type TImageTst  is array (0 to (8*17)-1) of std_logic_vector (31 downto 0);
constant C_TST_IMAGE : TImageTst:=(
--//Y0
(CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#041#, 8)&CONV_STD_LOGIC_VECTOR(10#034#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#045#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y1
(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#041#, 8)&CONV_STD_LOGIC_VECTOR(10#032#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#045#, 8)&CONV_STD_LOGIC_VECTOR(10#047#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y2
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#037#, 8)&CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#049#, 8)&CONV_STD_LOGIC_VECTOR(10#044#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y3
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#032#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#029#, 8)&CONV_STD_LOGIC_VECTOR(10#039#, 8)&CONV_STD_LOGIC_VECTOR(10#045#, 8)&CONV_STD_LOGIC_VECTOR(10#039#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y4
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#038#, 8)&CONV_STD_LOGIC_VECTOR(10#036#, 8)&CONV_STD_LOGIC_VECTOR(10#034#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y5
(CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#059#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#031#, 8)&CONV_STD_LOGIC_VECTOR(10#031#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#029#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y6
(CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#032#, 8)&CONV_STD_LOGIC_VECTOR(10#050#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y7
(CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y8
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#007#, 8)&CONV_STD_LOGIC_VECTOR(10#008#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y9
(CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y10
(CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y11
(CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#009#, 8)&CONV_STD_LOGIC_VECTOR(10#009#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y12
(CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y13
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y14
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y15
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)),  --//28..31


--//Y16
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8))  --//28..31

);

component vsobel_main
generic(
G_SIM : string:="OFF"
);
port
(
-------------------------------
-- ����������
-------------------------------
p_in_cfg_bypass            : in    std_logic;
p_in_cfg_pix_count         : in    std_logic_vector(15 downto 0);
p_in_cfg_row_count         : in    std_logic_vector(15 downto 0);
p_in_cfg_ctrl              : in    std_logic_vector(1 downto 0);

--//--------------------------
--//Upstream Port
--//--------------------------
p_in_upp_data              : in    std_logic_vector(31 downto 0);
p_in_upp_wd                : in    std_logic;
p_out_upp_rdy_n            : out   std_logic;

--//--------------------------
--//Downstream Port
--//--------------------------
p_in_dwnp_rdy_n            : in    std_logic;
p_out_dwnp_wd              : out   std_logic;
p_out_dwnp_data            : out   std_logic_vector(31 downto 0);

p_out_dwnp_dx              : out   std_logic_vector(7 downto 0);
p_out_dwnp_dy              : out   std_logic_vector(7 downto 0);
p_out_dwnp_grad            : out   std_logic_vector(7 downto 0);

-------------------------------
--���������������
-------------------------------
p_in_tst_ctrl              : in    std_logic_vector(31 downto 0);
p_out_tst                  : out   std_logic_vector(31 downto 0);

-------------------------------
--System
-------------------------------
p_in_clk            : in    std_logic;
p_in_rst            : in    std_logic
);
end component;

component vsobel_fifo
port (
din        : IN  std_logic_VECTOR(31 downto 0);
wr_en      : IN  std_logic;

dout       : OUT std_logic_VECTOR(31 downto 0);
rd_en      : IN  std_logic;

empty      : OUT std_logic;
full       : OUT std_logic;
almost_full: OUT std_logic;

clk        : IN  std_logic;
rst        : IN  std_logic
);
end component;


signal p_in_clk                       : std_logic := '0';
signal p_in_rst                       : std_logic := '0';

signal p_in_cfg_bypass                : std_logic;
--signal p_in_cfg_colorfst              : std_logic_vector(1 downto 0); --//0/1/2 - R/G/B
signal p_in_cfg_pix_count             : std_logic_vector(15 downto 0);
signal p_in_cfg_row_count             : std_logic_vector(15 downto 0);
signal p_in_cfg_ctrl                  : std_logic_vector(1 downto 0);

signal tst_data_out                   : std_logic_vector(31 downto 0);
signal p_in_upp_wd                    : std_logic;
signal p_out_upp_rdy_n                : std_logic;

signal p_out_dwnp_data                : std_logic_vector(31 downto 0);
signal p_out_dwnp_wd                  : std_logic;
signal p_in_dwnp_rdy_n                : std_logic;

signal i_fifoin_dout                  : std_logic_vector(31 downto 0);
signal i_fifoin_rd                    : std_logic;
signal i_fifoin_empty                 : std_logic;
signal i_fifoin_full                  : std_logic;

signal tst_mnl_vfr_count              : std_logic_vector(7 downto 0);
signal tst_mnl_pix_count              : std_logic_vector(15 downto 0);
signal tst_mnl_row_count              : std_logic_vector(15 downto 0);
signal tst_mnl_rowpuase_count         : std_logic_vector(15 downto 0);

signal tst_vfr_count                  : std_logic_vector(7 downto 0);
signal tst_puse_count                 : std_logic_vector(15 downto 0);
signal tst_row_count                  : std_logic_vector(15 downto 0);
signal tst_pix_count                  : std_logic_vector(15 downto 0);
signal tst_data                       : std_logic_vector(7 downto 0);
signal mnl_write_testdata             : std_logic;

signal tst_mnl_frpuase_count          : std_logic_vector(7 downto 0);
signal tst_frpuase_count              : std_logic_vector(7 downto 0);

signal mnl_use_gen_dwnp_rdy           : std_logic;
signal mnl_dwnp_rdy_n                 : std_logic;
signal i_dwnp_rdy_n                   : std_logic;

signal adr_image_out                  : std_logic_vector(7 downto 0);
signal tst_image_out                  : std_logic_vector(31 downto 0);

signal i_sobel_grad                   : std_logic_vector(7 downto 0);
signal tst_dwnp_pix                   : std_logic_vector(tst_mnl_pix_count'range);
signal tst_dwnp_row                   : std_logic_vector(31 downto 0);
signal tst_dwnp_count                 : std_logic_vector(31 downto 0);

--Main
begin



m_vsobel: vsobel_main
generic map(
G_SIM => "ON"
)
port map
(
-------------------------------
-- ����������
-------------------------------
p_in_cfg_bypass            => p_in_cfg_bypass,
p_in_cfg_pix_count         => p_in_cfg_pix_count,
p_in_cfg_row_count         => p_in_cfg_row_count,
p_in_cfg_ctrl              => p_in_cfg_ctrl,

--//--------------------------
--//Upstream Port
--//--------------------------
p_in_upp_data              => i_fifoin_dout,
p_in_upp_wd                => i_fifoin_rd,
p_out_upp_rdy_n            => p_out_upp_rdy_n,

--//--------------------------
--//Downstream Port
--//--------------------------
p_in_dwnp_rdy_n            => p_in_dwnp_rdy_n,
p_out_dwnp_wd              => p_out_dwnp_wd,
p_out_dwnp_data            => p_out_dwnp_data,

p_out_dwnp_dx              => open,
p_out_dwnp_dy              => open,
p_out_dwnp_grad            => i_sobel_grad,

-------------------------------
--���������������
-------------------------------
p_in_tst_ctrl              => "00000000000000000000000000000000",
p_out_tst                  => open,

-------------------------------
--System
-------------------------------
p_in_clk            => p_in_clk,
p_in_rst            => p_in_rst
);

m_fifo_in : vsobel_fifo
port map
(
din         => tst_image_out,--tst_data_out,
wr_en       => p_in_upp_wd,
--wr_clk      => p_in_upp_clk,

dout        => i_fifoin_dout,
rd_en       => i_fifoin_rd,
--rd_clk      => p_in_dwnp_clk,

empty       => i_fifoin_empty,
full        => open,
almost_full => i_fifoin_full,

clk         => p_in_clk,
rst         => p_in_rst
);

i_fifoin_rd<=not i_fifoin_empty and not p_out_upp_rdy_n;


clk_in_generator : process
begin
  p_in_clk<='0';
  wait for i_clk_period/2;
  p_in_clk<='1';
  wait for i_clk_period/2;
end process;


p_in_rst<='1','0' after 1 us;


--//----------------------------------------------------------
--//��������� ������������
--//----------------------------------------------------------
p_in_cfg_bypass<='0';--//0/1 - ���������� ������ �����/1 bypss

p_in_cfg_ctrl(0)<='0';-- 1/0 - ������ ������ ������������ ������� (dx^2 + dy^2)^0.5
p_in_cfg_ctrl(1)<='0';-- 1/0 - dx/2 � dy/2 /��� �������

--//������������� ��������� ��������� ������:
p_in_cfg_pix_count<=CONV_STD_LOGIC_VECTOR(10#06#, p_in_cfg_pix_count'length); --
p_in_cfg_row_count<=CONV_STD_LOGIC_VECTOR(10#16#, p_in_cfg_row_count'length); --
tst_mnl_vfr_count<=CONV_STD_LOGIC_VECTOR(16#01#, 8); --

tst_mnl_rowpuase_count<=CONV_STD_LOGIC_VECTOR(16#0F#, tst_mnl_rowpuase_count'length); --//����� ����� ��������
tst_mnl_frpuase_count<=CONV_STD_LOGIC_VECTOR(16#08#, tst_mnl_frpuase_count'length); --//����� ����� �������

--// 1/0 ������������/�� ������������� waveform ��� ������� p_in_dwnp_rdy_n
mnl_use_gen_dwnp_rdy<='0';




--//----------------------------------------------------------
--//
--//----------------------------------------------------------
p_in_dwnp_rdy_n<=i_dwnp_rdy_n when mnl_use_gen_dwnp_rdy='1' else '0';


tst_mnl_pix_count  <=p_in_cfg_pix_count;   --//���-�� ��������
tst_mnl_row_count  <=p_in_cfg_row_count;   --//���-�� �����

mnl_write_testdata<='0','1' after 2.5 us;


mnl_dwnp_rdy_n<='0',
                '1' after 2.5 us, '0' after 2.65654 us,
                '1' after 2.685 us, '1' after 2.6987 us,
                '1' after 2.8 us, '0' after 2.987 us,
                '1' after 3.0 us, '0' after 3.1234 us,
                '1' after 3.15 us, '0' after 3.18 us,
                '1' after 3.2 us, '0' after 3.23 us,
                '1' after 3.26 us, '0' after 3.3 us,
                '1' after 3.36 us,'0' after 3.39 us,
                '1' after 3.41 us,'0' after 3.43 us,
                '1' after 3.45 us,'0' after 3.46 us,
                '1' after 3.47 us,'0' after 3.48 us,
                '1' after 3.50 us,'0' after 3.51 us,
                '1' after 3.52 us,'0' after 3.5278 us,
                '1' after 3.53 us,'0' after 3.54 us,
                '1' after 3.55 us,'0' after 3.58 us,
                '1' after 3.63 us,'0' after 3.65 us,
                '1' after 3.70 us,'0' after 3.80 us,
                '1' after 3.84 us,'0' after 3.86 us,
                '1' after 3.89 us,'0' after 3.95 us,
                '1' after 4.0 us, '0' after 4.0678 us;


adr_image_out(7 downto 0)<=tst_row_count(4 downto 0)&tst_pix_count(2 downto 0);
tst_image_out<=C_TST_IMAGE(CONV_INTEGER(adr_image_out));

--//��������� �������� ������
process(p_in_rst,p_in_clk)
  variable GUI_line : LINE;--������ ��_ ������ � ModelSim
begin
  if p_in_rst='1' then
    tst_vfr_count<=(others=>'0');
    tst_row_count<=(others=>'0');
    tst_puse_count<=(others=>'0');
    tst_pix_count<=(others=>'0');
    tst_frpuase_count<=(others=>'0');
    tst_data<=CONV_STD_LOGIC_VECTOR(16#2#, tst_data'length); --//
    tst_data_out<=(others=>'0');
    p_in_upp_wd<='0';
    i_dwnp_rdy_n<='0';

  elsif p_in_clk'event and p_in_clk='1' then
    i_dwnp_rdy_n<=mnl_dwnp_rdy_n;

    if mnl_write_testdata='1' then

--      if p_out_upp_rdy_n='0' then
      if i_fifoin_full='0' then

        if tst_pix_count=tst_mnl_pix_count-1 then
          if tst_row_count=tst_mnl_row_count-1 then
            if tst_vfr_count=tst_mnl_vfr_count-1 then
              tst_row_count<=tst_row_count;
              tst_pix_count<=tst_pix_count;
              tst_vfr_count<=tst_vfr_count;
            else
              if tst_frpuase_count=tst_mnl_frpuase_count then
                tst_frpuase_count<=(others=>'0');
                tst_row_count<=(others=>'0');
                tst_pix_count<=(others=>'0');
                tst_vfr_count<=tst_vfr_count+1;
              else
                tst_frpuase_count<=tst_frpuase_count+1;
              end if;
            end if;
            p_in_upp_wd<='0';
          else
            if tst_puse_count=tst_mnl_rowpuase_count then
              tst_puse_count<=(others=>'0');

              tst_row_count<=tst_row_count+1;
              tst_pix_count<=(others=>'0');
              p_in_upp_wd<='1';

              tst_data<=tst_data+8;
              tst_data_out(7 downto 0)  <=tst_data;
              tst_data_out(15 downto 8) <=tst_data+2;
              tst_data_out(23 downto 16)<=tst_data+4;
              tst_data_out(31 downto 24)<=tst_data+6;

            else
              p_in_upp_wd<='0';
              tst_puse_count<=tst_puse_count+1;
            end if;
          end if;

        else
          if p_in_upp_wd='1' then
          tst_pix_count<=tst_pix_count+1;
          end if;
          p_in_upp_wd<='1';

--          tst_data<=tst_data+4;
--          tst_data_out(7 downto 0)  <=tst_data;
--          tst_data_out(15 downto 8) <=tst_data+1;
--          tst_data_out(23 downto 16)<=tst_data+2;
--          tst_data_out(31 downto 24)<=tst_data+3;

          tst_data<=tst_data+8;
          tst_data_out(7 downto 0)  <=tst_data;
          tst_data_out(15 downto 8) <=tst_data+2;
          tst_data_out(23 downto 16)<=tst_data+4;
          tst_data_out(31 downto 24)<=tst_data+6;

        end if;
      else
        p_in_upp_wd<='0';
      end if;
    else
      p_in_upp_wd<='0';
    end if;

  end if;
end process;


--//������� � ������� ModelSim ��������� ���������� ��������� �������
process(p_in_rst,p_in_clk)
  variable GUI_line : LINE;--������ ��_ ������ � ModelSim
begin
  if p_in_rst='1' then
    tst_dwnp_pix<=(others=>'0');
    tst_dwnp_row<=(others=>'0');
  elsif p_in_clk'event and p_in_clk='1' then

    if p_out_dwnp_wd='1' and p_in_dwnp_rdy_n='0' then
        if tst_dwnp_pix=(tst_dwnp_pix'range=>'0') then
          write(GUI_line, string'("Result: Line("));
          write(GUI_line, itoa(CONV_INTEGER(tst_dwnp_row)));--//������ ����� � DEC
          write(GUI_line, string'(") "));
        end if;

        write(GUI_line, itoa(CONV_INTEGER(i_sobel_grad)));--//������ ����� � DEC
        write(GUI_line, string'(","));

        if tst_dwnp_pix=((tst_mnl_pix_count(13 downto 0)&"00")-1) then
          tst_dwnp_pix<=(others=>'0');
          tst_dwnp_row<=tst_dwnp_row+1;
          writeline(output, GUI_line);--������� ������ GUI_line � ModelSim
        else
          tst_dwnp_pix<=tst_dwnp_pix+1;
        end if;
    end if;

  end if;
end process;

--process(p_in_rst,p_in_clk)
--  variable GUI_line : LINE;--������ ��_ ������ � ModelSim
--begin
--  if p_in_rst='1' then
--    tst_dwnp_count<=(others=>'0');
--  elsif p_in_clk'event and p_in_clk='1' then
--
--    if p_out_dwnp_wd='1' and p_in_dwnp_rdy_n='0' then
--        tst_dwnp_count<=tst_dwnp_count+1;
--
--        write(GUI_line, string'("Result 2DW ("));
--        hwrite(GUI_line, tst_dwnp_count);--//������ ����� � HEX
--        write(GUI_line, string'(") : 0x"));
--        hwrite(GUI_line, p_out_dwnp_data);--//������ ����� � HEX
--        writeline(output, GUI_line);--������� ������ GUI_line � ModelSim
--    end if;
--
--  end if;
--end process;

--End Main
end;
