-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 26.10.2012 13:05:53
-- Module Name : eth_bram_prm
--
-- ����������/�������� :
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

entity eth_bram_prm is
port(
p_out_cfg_adr      : out  std_logic_vector(7 downto 0);
p_out_cfg_adr_ld   : out  std_logic;
p_out_cfg_adr_fifo : out  std_logic;

p_out_cfg_txdata   : out  std_logic_vector(15 downto 0);
p_out_cfg_wr       : out  std_logic;

p_in_clk  : in  std_logic;
p_in_rst  : in  std_logic
);
end eth_bram_prm;

architecture behavioral of eth_bram_prm is

constant CI_ETH_REG_CTRL : integer := 0;

signal i_addra : std_logic_vector(15 downto 0);
signal i_douta : std_logic_vector(31 downto 0);

type TEth_cfg_fsm is (
S_CFG_ETH_START,
S_CFG_ETH_MAC_DST0,
S_CFG_ETH_MAC_DST1,
S_CFG_ETH_MAC_DST2,
S_CFG_ETH_MAC_SRC0,
S_CFG_ETH_MAC_SRC1,
S_CFG_ETH_MAC_SRC2,
S_CFG_ETH_IP_DST0,
S_CFG_ETH_IP_DST1,
S_CFG_ETH_IP_SRC0,
S_CFG_ETH_IP_SRC1,
S_CFG_ETH_PORT_DST,
S_CFG_ETH_PORT_SRC,
S_CFG_ETH_CTRL,
S_CFG_ETH_DONE
);
signal fsm_ethcfg_cs: TEth_cfg_fsm;

signal i_eth_prm_a   : std_logic_vector(4 downto 0);
signal i_eth_prm_d   : std_logic_vector(15 downto 0);

signal i_eth_cfg_radr                  : std_logic_vector(7 downto 0);
signal i_eth_cfg_radr_ld               : std_logic;
signal i_eth_cfg_radr_fifo             : std_logic;
signal i_eth_cfg_wr                    : std_logic;
signal i_eth_cfg_txd                   : std_logic_vector(15 downto 0);


--MAIN
begin


p_out_cfg_adr      <= i_eth_cfg_radr;
p_out_cfg_adr_ld   <= i_eth_cfg_radr_ld;
p_out_cfg_adr_fifo <= i_eth_cfg_radr_fifo;

p_out_cfg_txdata   <= i_eth_cfg_txd;
p_out_cfg_wr       <= i_eth_cfg_wr;

process(p_in_rst,p_in_clk)
begin
  if p_in_rst = '1' then
    i_eth_prm_a <= (others=>'0');
  elsif rising_edge(p_in_clk) then
    if fsm_ethcfg_cs /= S_CFG_ETH_DONE then --and p_in_clk.rdy='1' then
      i_eth_prm_a <= i_eth_prm_a + 1;
    else
      i_eth_prm_a <= (others=>'0');
    end if;
  end if;
end process;

process(p_in_rst,p_in_clk)
begin
  if p_in_rst = '1' then
    fsm_ethcfg_cs<=S_CFG_ETH_START;

    i_eth_cfg_radr<=(others=>'0');
    i_eth_cfg_radr_ld<='0';
    i_eth_cfg_radr_fifo<='0';

    i_eth_cfg_txd<=(others=>'0');
    i_eth_cfg_wr<='0';
--    i_eth_cfg_done<='0';

  elsif rising_edge(p_in_clk) then

    case fsm_ethcfg_cs is

      --
      when S_CFG_ETH_START =>

--        if p_in_rdy='1' then
        i_eth_cfg_radr_ld<='1';
        i_eth_cfg_radr_fifo<='0';
        i_eth_cfg_wr<='0';
        i_eth_cfg_radr<=CONV_STD_LOGIC_VECTOR(CI_ETH_REG_CTRL, i_eth_cfg_radr'length);
        fsm_ethcfg_cs<=S_CFG_ETH_CTRL;
--        end if;

      --Set CTRL
      when S_CFG_ETH_CTRL =>
        i_eth_cfg_radr_ld<='0';
        i_eth_cfg_radr_fifo<='0';
        i_eth_cfg_wr<='1';
        i_eth_cfg_txd(8*2-1 downto 8*0)<=i_eth_prm_d(8*2-1 downto 8*0);
        fsm_ethcfg_cs<=S_CFG_ETH_MAC_DST0;

      --Set MAC/DST
      when S_CFG_ETH_MAC_DST0 =>
        i_eth_cfg_radr_ld<='0';
        i_eth_cfg_radr_fifo<='0';
        i_eth_cfg_wr<='1';
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_MAC_DST1;

      when S_CFG_ETH_MAC_DST1 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_MAC_DST2;

      when S_CFG_ETH_MAC_DST2 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_MAC_SRC0;

      --Set MAC/SRC
      when S_CFG_ETH_MAC_SRC0 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_MAC_SRC1;

      when S_CFG_ETH_MAC_SRC1 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_MAC_SRC2;

      when S_CFG_ETH_MAC_SRC2 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_IP_DST0;

      --Set IP/DST
      when S_CFG_ETH_IP_DST0 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_IP_DST1;

      when S_CFG_ETH_IP_DST1 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_IP_SRC0;

      --Set IP/SRC
      when S_CFG_ETH_IP_SRC0 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_IP_SRC1;

      when S_CFG_ETH_IP_SRC1 =>
        i_eth_cfg_txd(8*1-1 downto 8*0)<=i_eth_prm_d(8*1-1 downto 8*0);
        i_eth_cfg_txd(8*2-1 downto 8*1)<=i_eth_prm_d(8*2-1 downto 8*1);
        fsm_ethcfg_cs<=S_CFG_ETH_PORT_DST;

      --Set PORT/DST
      when S_CFG_ETH_PORT_DST =>
        i_eth_cfg_txd(8*2-1 downto 8*0)<=i_eth_prm_d(8*2-1 downto 8*0);
        fsm_ethcfg_cs<=S_CFG_ETH_PORT_SRC;

      --Set PORT/SRC
      when S_CFG_ETH_PORT_SRC =>
        i_eth_cfg_txd(8*2-1 downto 8*0)<=i_eth_prm_d(8*2-1 downto 8*0);
        fsm_ethcfg_cs<=S_CFG_ETH_DONE;

      when S_CFG_ETH_DONE =>
        i_eth_cfg_wr<='0';
--        i_eth_cfg_done<='1';

    end case;
  end if;
end process;


   m_core : RAMB36
   generic map (
      DOA_REG => 0,  -- Optional output register on A port (0 or 1)
      DOB_REG => 0,  -- Optional output register on B port (0 or 1)
      INIT_A => X"000000000", -- Initial values on A output port
      INIT_B => X"000000000", -- Initial values on B output port
      RAM_EXTENSION_A => "NONE",  -- "UPPER", "LOWER" or "NONE" when cascaded
      RAM_EXTENSION_B => "NONE",  -- "UPPER", "LOWER" or "NONE" when cascaded
      READ_WIDTH_A => 18,   -- Valid values are 1, 2, 4, 9, 18, or 36
      READ_WIDTH_B => 18,   -- Valid values are 1, 2, 4, 9, 18, or 36
      SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY",
                                    -- "GENERATE_X_ONLY" or "NONE"
      SIM_MODE => "SAFE", -- Simulation: "SAFE" vs "FAST", see "Synthesis and Simulation
                          -- Design Guide" for details
      SRVAL_A => X"000000000",   -- Set/Reset value for A port output
      SRVAL_B => X"000000000",   -- Set/Reset value for B port output
      WRITE_MODE_A => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
      WRITE_MODE_B => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
      WRITE_WIDTH_A => 18,  -- Valid values are 1, 2, 3, 4, 9, 18, 36
      WRITE_WIDTH_B => 18,  -- Valid values are 1, 2, 3, 4, 9, 18, 36
      -- The following INIT_xx declarations specify the initial contents of the RAM
      INIT_00 => X"0000000000000BB80BB8EB07010A7D07010A000000DC0800DA31CEBAE6900000", --default : DHCP-on; FPGA mac/ip/port - 00:08:DC:00:00/10.1.7.235/3000; HOST mac/ip/port - 90:E6:BA:CE:31:DA/10.1.7.125/3000
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      CASCADEOUTLATA => open,--CASCADEOUTLATA,   -- 1-bit cascade A latch output
      CASCADEOUTLATB => open,--CASCADEOUTLATB,   -- 1-bit cascade B latch output
      CASCADEOUTREGA => open,--CASCADEOUTREGA,   -- 1-bit cascade A register output
      CASCADEOUTREGB => open,--CASCADEOUTREGB,   -- 1-bit cascade B register output
      DOA => i_douta, -- 32-bit A port data output
      DOB => open, -- 32-bit B port data output
      DOPA => open,  -- 4-bit A port parity data output
      DOPB => open,  -- 4-bit B port parity data output
      ADDRA => i_addra, -- 16-bit A port address input
      ADDRB => (others=>'0'), -- 16-bit B port address input
      CASCADEINLATA => '0',--CASCADEINLATA,  -- 1-bit cascade A latch input
      CASCADEINLATB => '0',--CASCADEINLATB,  -- 1-bit cascade B latch input
      CASCADEINREGA => '0',--CASCADEINREGA,  -- 1-bit cascade A register input
      CASCADEINREGB => '0',--CASCADEINREGB,  -- 1-bit cascade B register input
      CLKA => p_in_clk,  -- 1-bit A port clock input
      CLKB => p_in_clk,  -- 1 bit B port clock input
      DIA => (others=>'0'), -- 32-bit A port data input
      DIB => (others=>'0'), -- 32-bit B port data input
      DIPA => (others=>'0'),  -- 4-bit A port parity data input
      DIPB => (others=>'0'),  -- 4-bit B port parity data input
      ENA => '1', -- 1-bit A port enable input
      ENB => '1', -- 1-bit B port enable input
      REGCEA => '0', -- 1-bit A port register enable input
      REGCEB => '0', -- 1-bit B port register enable input
      SSRA => '0',  -- 1-bit A port set/reset input
      SSRB => '0',  -- 1-bit B port set/reset input
      WEA => (others=>'0'), -- 4-bit A port write enable input
      WEB => (others=>'0')  -- 4-bit B port write enable input
   );

i_addra <= '0' & "000000" & i_eth_prm_a(4 downto 0) & "0000";

gen : for i in 0 to 15 generate
i_eth_prm_d(i) <= i_douta(i);
end generate gen;

--END MAIN
end behavioral;

