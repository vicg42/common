//-----------------------------------------------------------------------
// author    : Golovachenko Victor
//------------------------------------------------------------------------

module filter_median_7x7 #(
    parameter LINE_SIZE_MAX = 1024,
    parameter PIXEL_WIDTH = 12
)(
    input bypass,

    //input resolution X * Y
    input [PIXEL_WIDTH-1:0] di_i,
    input                   de_i,
    input                   hs_i,
    input                   vs_i,

    //output resolution (X - 4) * (Y - 4)
    output [PIXEL_WIDTH-1:0] do_o, //
    output                   de_o, //
    output                   hs_o, //
    output                   vs_o, //

    output [PIXEL_WIDTH-1:0] bypass_o, //

    input clk,
    input rst
);

function [PIXEL_WIDTH*2-1:0] Sort2;
    input [PIXEL_WIDTH-1:0] x1;
    input [PIXEL_WIDTH-1:0] x2;
    if (x1 > x2)
        Sort2 = {x2, x1};
    else
        Sort2 = {x1, x2};
endfunction


localparam KERNEL_SIZE = 49;

wire [(PIXEL_WIDTH*KERNEL_SIZE)-1:0] xi;
wire [(PIXEL_WIDTH*KERNEL_SIZE)-1:0] xo;

reg [PIXEL_WIDTH-1:0] s00 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s01 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s02 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s03 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s04 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s05 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s06 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s07 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s08 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s09 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s10 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s11 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s12 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s13 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s14 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s15 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s16 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s17 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s18 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s19 [(KERNEL_SIZE)-1:0];
reg [PIXEL_WIDTH-1:0] s20 [(KERNEL_SIZE)-1:0];

wire de;
wire hs;
wire vs;
reg [0:20] sr_de = 0;
reg [0:20] sr_hs = 0;
reg [0:20] sr_vs = 0;
reg [PIXEL_WIDTH-1:0] sr_bypass_data [0:20];

filter_core_7x7 #(
    .DE_I_PERIOD(0),
    .LINE_SIZE_MAX (LINE_SIZE_MAX),
    .DATA_WIDTH (PIXEL_WIDTH)
) filter_core_7x7 (
    .bypass(1'b0),

    .di_i(di_i),
    .de_i(de_i),
    .hs_i(hs_i),
    .vs_i(vs_i),

    //output resolution (X - 6) * (Y - 6)
    //pixel pattern:
    //line[0]: x00 x01 x02 x03 x04 x05 x06
    //line[1]: x07 x08 x09 x10 x11 x12 x13
    //line[2]: x14 x15 x16 x17 x18 x19 x20
    //line[3]: x21 x22 x23 x24 x25 x26 x27
    //line[4]: x28 x29 x30 x31 x32 x33 x34
    //line[5]: x35 x36 x37 x38 x39 x40 x41
    //line[6]: x42 x43 x44 x45 x46 x47 x48
    .x00(xi[(PIXEL_WIDTH*( 0)) +: PIXEL_WIDTH]),
    .x01(xi[(PIXEL_WIDTH*( 1)) +: PIXEL_WIDTH]),
    .x02(xi[(PIXEL_WIDTH*( 2)) +: PIXEL_WIDTH]),
    .x03(xi[(PIXEL_WIDTH*( 3)) +: PIXEL_WIDTH]),
    .x04(xi[(PIXEL_WIDTH*( 4)) +: PIXEL_WIDTH]),
    .x05(xi[(PIXEL_WIDTH*( 5)) +: PIXEL_WIDTH]),
    .x06(xi[(PIXEL_WIDTH*( 6)) +: PIXEL_WIDTH]),
    .x07(xi[(PIXEL_WIDTH*( 7)) +: PIXEL_WIDTH]),
    .x08(xi[(PIXEL_WIDTH*( 8)) +: PIXEL_WIDTH]),
    .x09(xi[(PIXEL_WIDTH*( 9)) +: PIXEL_WIDTH]),
    .x10(xi[(PIXEL_WIDTH*(10)) +: PIXEL_WIDTH]),
    .x11(xi[(PIXEL_WIDTH*(11)) +: PIXEL_WIDTH]),
    .x12(xi[(PIXEL_WIDTH*(12)) +: PIXEL_WIDTH]),
    .x13(xi[(PIXEL_WIDTH*(13)) +: PIXEL_WIDTH]),
    .x14(xi[(PIXEL_WIDTH*(14)) +: PIXEL_WIDTH]),
    .x15(xi[(PIXEL_WIDTH*(15)) +: PIXEL_WIDTH]),
    .x16(xi[(PIXEL_WIDTH*(16)) +: PIXEL_WIDTH]),
    .x17(xi[(PIXEL_WIDTH*(17)) +: PIXEL_WIDTH]),
    .x18(xi[(PIXEL_WIDTH*(18)) +: PIXEL_WIDTH]),
    .x19(xi[(PIXEL_WIDTH*(19)) +: PIXEL_WIDTH]),
    .x20(xi[(PIXEL_WIDTH*(20)) +: PIXEL_WIDTH]),
    .x21(xi[(PIXEL_WIDTH*(21)) +: PIXEL_WIDTH]),
    .x22(xi[(PIXEL_WIDTH*(22)) +: PIXEL_WIDTH]),
    .x23(xi[(PIXEL_WIDTH*(23)) +: PIXEL_WIDTH]),
    .x24(xi[(PIXEL_WIDTH*(24)) +: PIXEL_WIDTH]),
    .x25(xi[(PIXEL_WIDTH*(25)) +: PIXEL_WIDTH]),
    .x26(xi[(PIXEL_WIDTH*(26)) +: PIXEL_WIDTH]),
    .x27(xi[(PIXEL_WIDTH*(27)) +: PIXEL_WIDTH]),
    .x28(xi[(PIXEL_WIDTH*(28)) +: PIXEL_WIDTH]),
    .x29(xi[(PIXEL_WIDTH*(29)) +: PIXEL_WIDTH]),
    .x30(xi[(PIXEL_WIDTH*(30)) +: PIXEL_WIDTH]),
    .x31(xi[(PIXEL_WIDTH*(31)) +: PIXEL_WIDTH]),
    .x32(xi[(PIXEL_WIDTH*(32)) +: PIXEL_WIDTH]),
    .x33(xi[(PIXEL_WIDTH*(33)) +: PIXEL_WIDTH]),
    .x34(xi[(PIXEL_WIDTH*(34)) +: PIXEL_WIDTH]),
    .x35(xi[(PIXEL_WIDTH*(35)) +: PIXEL_WIDTH]),
    .x36(xi[(PIXEL_WIDTH*(36)) +: PIXEL_WIDTH]),
    .x37(xi[(PIXEL_WIDTH*(37)) +: PIXEL_WIDTH]),
    .x38(xi[(PIXEL_WIDTH*(38)) +: PIXEL_WIDTH]),
    .x39(xi[(PIXEL_WIDTH*(39)) +: PIXEL_WIDTH]),
    .x40(xi[(PIXEL_WIDTH*(40)) +: PIXEL_WIDTH]),
    .x41(xi[(PIXEL_WIDTH*(41)) +: PIXEL_WIDTH]),
    .x42(xi[(PIXEL_WIDTH*(42)) +: PIXEL_WIDTH]),
    .x43(xi[(PIXEL_WIDTH*(43)) +: PIXEL_WIDTH]),
    .x44(xi[(PIXEL_WIDTH*(44)) +: PIXEL_WIDTH]),
    .x45(xi[(PIXEL_WIDTH*(45)) +: PIXEL_WIDTH]),
    .x46(xi[(PIXEL_WIDTH*(46)) +: PIXEL_WIDTH]),
    .x47(xi[(PIXEL_WIDTH*(47)) +: PIXEL_WIDTH]),
    .x48(xi[(PIXEL_WIDTH*(48)) +: PIXEL_WIDTH]),

    .de_o(de),
    .hs_o(hs),
    .vs_o(vs),

    .clk (clk),
    .rst (rst)
);

// -------------------------------------------------------------------------
// pixel buffer, making following pixel pattern:
// -------------------------------------------------------------------------
// x00 x01 x02 x03 x04 x05 x06
// x07 x08 x09 x10 x11 x12 x13
// x14 x15 x16 x17 x18 x19 x20
// x21 x22 x23 x24 x25 x26 x27
// x28 x29 x30 x31 x32 x33 x34
// x35 x36 x37 x38 x39 x40 x41
// x42 x43 x44 x45 x46 x47 x48



integer a,a1,b,b1,c,c1,d,d1,e;
always @(posedge clk) begin
    //stage0
    for (a=0; a<32; a=a+2) begin
        {s00[(a+0)], s00[(a+1)]} <= Sort2(xi[(PIXEL_WIDTH*(a+0)) +: PIXEL_WIDTH], xi[(PIXEL_WIDTH*(a+1)) +: PIXEL_WIDTH]);
    end
    for (a1=32; a1<48; a1=a1+2) begin
        {s00[(a1+0)], s00[(a1+1)]} <= Sort2(xi[(PIXEL_WIDTH*(a1+0)) +: PIXEL_WIDTH], xi[(PIXEL_WIDTH*(a1+1)) +: PIXEL_WIDTH]);
    end
    s00[(48)] <= xi[(PIXEL_WIDTH*(48)) +: PIXEL_WIDTH];

    sr_bypass_data[0] <= xi[(PIXEL_WIDTH*(24)) +: PIXEL_WIDTH];
    sr_de[0] <= de;
    sr_hs[0] <= hs;
    sr_vs[0] <= vs;

    for (b=0; b<32; b=b+4) begin
        //stage1
        {s01[(b+0)], s01[(b+2)]} <= Sort2(s00[(b+0)], s00[(b+2)]);
        {s01[(b+1)], s01[(b+3)]} <= Sort2(s00[(b+1)], s00[(b+3)]);

        //stage2
                    s02[(b+0)] <= s01[(b+0)];
        {s02[(b+1)], s02[(b+2)]} <= Sort2(s01[(b+1)], s01[(b+2)]);
                    s02[(b+3)] <= s01[(b+3)];
    end
    for (b1=32; b1<48; b1=b1+4) begin
        //stage1
        {s01[(b1+0)], s01[(b1+2)]} <= Sort2(s00[(b1+0)], s00[(b1+2)]);
        {s01[(b1+1)], s01[(b1+3)]} <= Sort2(s00[(b1+1)], s00[(b1+3)]);

        //stage2
                    s02[(b1+0)] <= s01[(b1+0)];
        {s02[(b1+1)], s02[(b1+2)]} <= Sort2(s01[(b1+1)], s01[(b1+2)]);
                    s02[(b1+3)] <= s01[(b1+3)];
    end
    s01[(48)] <= s00[(48)];
    s02[(48)] <= s01[(48)];
    sr_bypass_data[1] <= sr_bypass_data[0];
    sr_de[1] <= sr_de[0];
    sr_hs[1] <= sr_hs[0];
    sr_vs[1] <= sr_vs[0];
    sr_bypass_data[2] <= sr_bypass_data[1];
    sr_de[2] <= sr_de[1];
    sr_hs[2] <= sr_hs[1];
    sr_vs[2] <= sr_vs[1];


    for (c=0; c<32; c=c+8) begin
        //stage3
        {s03[(c+0)], s03[(c+4)]} <= Sort2(s02[(c+0)], s02[(c+4)]);
        {s03[(c+1)], s03[(c+5)]} <= Sort2(s02[(c+1)], s02[(c+5)]);
        {s03[(c+2)], s03[(c+6)]} <= Sort2(s02[(c+2)], s02[(c+6)]);
        {s03[(c+3)], s03[(c+7)]} <= Sort2(s02[(c+3)], s02[(c+7)]);

        //stage4
                    s04[(c+0)] <= s03[(c+0)];
                    s04[(c+1)] <= s03[(c+1)];
        {s04[(c+2)], s04[(c+4)]} <= Sort2(s03[(c+2)], s03[(c+4)]);
        {s04[(c+3)], s04[(c+5)]} <= Sort2(s03[(c+3)], s03[(c+5)]);
                    s04[(c+6)] <= s03[(c+6)];
                    s04[(c+7)] <= s03[(c+7)];

        //stage5
                    s05[(c+0)] <= s04[(c+0)];
        {s05[(c+1)], s05[(c+2)]} <= Sort2(s04[(c+1)], s04[(c+2)]);
        {s05[(c+3)], s05[(c+4)]} <= Sort2(s04[(c+3)], s04[(c+4)]);
        {s05[(c+5)], s05[(c+6)]} <= Sort2(s04[(c+5)], s04[(c+6)]);
                    s05[(c+7)] <= s04[(c+7)];
    end
    for (c1=32; c1<48; c1=c1+8) begin
        //stage3
        {s03[(c1+0)], s03[(c1+4)]} <= Sort2(s02[(c1+0)], s02[(c1+4)]);
        {s03[(c1+1)], s03[(c1+5)]} <= Sort2(s02[(c1+1)], s02[(c1+5)]);
        {s03[(c1+2)], s03[(c1+6)]} <= Sort2(s02[(c1+2)], s02[(c1+6)]);
        {s03[(c1+3)], s03[(c1+7)]} <= Sort2(s02[(c1+3)], s02[(c1+7)]);

        //stage4
                    s04[(c1+0)] <= s03[(c1+0)];
                    s04[(c1+1)] <= s03[(c1+1)];
        {s04[(c1+2)], s04[(c1+4)]} <= Sort2(s03[(c1+2)], s03[(c1+4)]);
        {s04[(c1+3)], s04[(c1+5)]} <= Sort2(s03[(c1+3)], s03[(c1+5)]);
                    s04[(c1+6)] <= s03[(c1+6)];
                    s04[(c1+7)] <= s03[(c1+7)];

        //stage5
                    s05[(c1+0)] <= s04[(c1+0)];
        {s05[(c1+1)], s05[(c1+2)]} <= Sort2(s04[(c1+1)], s04[(c1+2)]);
        {s05[(c1+3)], s05[(c1+4)]} <= Sort2(s04[(c1+3)], s04[(c1+4)]);
        {s05[(c1+5)], s05[(c1+6)]} <= Sort2(s04[(c1+5)], s04[(c1+6)]);
                    s05[(c1+7)] <= s04[(c1+7)];
    end
    s03[(48)] <= s02[(48)];
    s04[(48)] <= s03[(48)];
    s05[(48)] <= s04[(48)];

    sr_bypass_data[3] <= sr_bypass_data[2];
    sr_de[3] <= sr_de[2];
    sr_hs[3] <= sr_hs[2];
    sr_vs[3] <= sr_vs[2];

    sr_bypass_data[4] <= sr_bypass_data[3];
    sr_de[4] <= sr_de[3];
    sr_hs[4] <= sr_hs[3];
    sr_vs[4] <= sr_vs[3];

    sr_bypass_data[5] <= sr_bypass_data[4];
    sr_de[5] <= sr_de[4];
    sr_hs[5] <= sr_hs[4];
    sr_vs[5] <= sr_vs[4];

    for (d=0; d<32; d=d+16) begin
        //stage6
        {s06[(d+0)], s06[(d+ 8)]} <= Sort2(s05[(d+0)], s05[(d+ 8)]);
        {s06[(d+1)], s06[(d+ 9)]} <= Sort2(s05[(d+1)], s05[(d+ 9)]);
        {s06[(d+2)], s06[(d+10)]} <= Sort2(s05[(d+2)], s05[(d+10)]);
        {s06[(d+3)], s06[(d+11)]} <= Sort2(s05[(d+3)], s05[(d+11)]);
        {s06[(d+4)], s06[(d+12)]} <= Sort2(s05[(d+4)], s05[(d+12)]);
        {s06[(d+5)], s06[(d+13)]} <= Sort2(s05[(d+5)], s05[(d+13)]);
        {s06[(d+6)], s06[(d+14)]} <= Sort2(s05[(d+6)], s05[(d+14)]);
        {s06[(d+7)], s06[(d+15)]} <= Sort2(s05[(d+7)], s05[(d+15)]);

        //stage7
                    s07[(d+0)] <= s06[(d+0)];
                    s07[(d+1)] <= s06[(d+1)];
                    s07[(d+2)] <= s06[(d+2)];
                    s07[(d+3)] <= s06[(d+3)];
        {s07[(d+4)], s07[(d+ 8)]} <= Sort2(s06[(d+4)], s06[(d+ 8)]);
        {s07[(d+5)], s07[(d+ 9)]} <= Sort2(s06[(d+5)], s06[(d+ 9)]);
        {s07[(d+6)], s07[(d+10)]} <= Sort2(s06[(d+6)], s06[(d+10)]);
        {s07[(d+7)], s07[(d+11)]} <= Sort2(s06[(d+7)], s06[(d+11)]);
                    s07[(d+12)] <= s06[(d+12)];
                    s07[(d+13)] <= s06[(d+13)];
                    s07[(d+14)] <= s06[(d+14)];
                    s07[(d+15)] <= s06[(d+15)];

        //stage8
                    s08[(d+0)] <= s07[(d+0)];
                    s08[(d+1)] <= s07[(d+1)];
        {s08[(d+ 2)], s08[(d+ 4)]} <= Sort2(s07[(d+ 2)], s07[(d+ 4)]);
        {s08[(d+ 3)], s08[(d+ 5)]} <= Sort2(s07[(d+ 3)], s07[(d+ 5)]);
        {s08[(d+ 6)], s08[(d+ 8)]} <= Sort2(s07[(d+ 6)], s07[(d+ 8)]);
        {s08[(d+ 7)], s08[(d+ 9)]} <= Sort2(s07[(d+ 7)], s07[(d+ 9)]);
        {s08[(d+10)], s08[(d+12)]} <= Sort2(s07[(d+10)], s07[(d+12)]);
        {s08[(d+11)], s08[(d+13)]} <= Sort2(s07[(d+11)], s07[(d+13)]);
                    s08[(d+14)] <= s07[(d+14)];
                    s08[(d+15)] <= s07[(d+15)];

        //stage9
                    s09[(d+0)] <= s08[(d+0)];
        {s09[(d+ 1)], s09[(d+ 2)]} <= Sort2(s08[(d+ 1)], s08[(d+ 2)]);
        {s09[(d+ 3)], s09[(d+ 4)]} <= Sort2(s08[(d+ 3)], s08[(d+ 4)]);
        {s09[(d+ 5)], s09[(d+ 6)]} <= Sort2(s08[(d+ 5)], s08[(d+ 6)]);
        {s09[(d+ 7)], s09[(d+ 8)]} <= Sort2(s08[(d+ 7)], s08[(d+ 8)]);
        {s09[(d+ 9)], s09[(d+10)]} <= Sort2(s08[(d+ 9)], s08[(d+10)]);
        {s09[(d+11)], s09[(d+12)]} <= Sort2(s08[(d+11)], s08[(d+12)]);
        {s09[(d+13)], s09[(d+14)]} <= Sort2(s08[(d+13)], s08[(d+14)]);
                    s09[(d+15)] <= s08[(d+15)];
    end
    for (d1=32; d1<48; d1=d1+16) begin
        //stage6
        {s06[(d1+0)], s06[(d1+ 8)]} <= Sort2(s05[(d1+0)], s05[(d1+ 8)]);
        {s06[(d1+1)], s06[(d1+ 9)]} <= Sort2(s05[(d1+1)], s05[(d1+ 9)]);
        {s06[(d1+2)], s06[(d1+10)]} <= Sort2(s05[(d1+2)], s05[(d1+10)]);
        {s06[(d1+3)], s06[(d1+11)]} <= Sort2(s05[(d1+3)], s05[(d1+11)]);
        {s06[(d1+4)], s06[(d1+12)]} <= Sort2(s05[(d1+4)], s05[(d1+12)]);
        {s06[(d1+5)], s06[(d1+13)]} <= Sort2(s05[(d1+5)], s05[(d1+13)]);
        {s06[(d1+6)], s06[(d1+14)]} <= Sort2(s05[(d1+6)], s05[(d1+14)]);
        {s06[(d1+7)], s06[(d1+15)]} <= Sort2(s05[(d1+7)], s05[(d1+15)]);

        //stage7
                    s07[(d1+0)] <= s06[(d1+0)];
                    s07[(d1+1)] <= s06[(d1+1)];
                    s07[(d1+2)] <= s06[(d1+2)];
                    s07[(d1+3)] <= s06[(d1+3)];
        {s07[(d1+4)], s07[(d1+ 8)]} <= Sort2(s06[(d1+4)], s06[(d1+ 8)]);
        {s07[(d1+5)], s07[(d1+ 9)]} <= Sort2(s06[(d1+5)], s06[(d1+ 9)]);
        {s07[(d1+6)], s07[(d1+10)]} <= Sort2(s06[(d1+6)], s06[(d1+10)]);
        {s07[(d1+7)], s07[(d1+11)]} <= Sort2(s06[(d1+7)], s06[(d1+11)]);
                    s07[(d1+12)] <= s06[(d1+12)];
                    s07[(d1+13)] <= s06[(d1+13)];
                    s07[(d1+14)] <= s06[(d1+14)];
                    s07[(d1+15)] <= s06[(d1+15)];

        //stage8
                    s08[(d1+0)] <= s07[(d1+0)];
                    s08[(d1+1)] <= s07[(d1+1)];
        {s08[(d1+ 2)], s08[(d1+ 4)]} <= Sort2(s07[(d1+ 2)], s07[(d1+ 4)]);
        {s08[(d1+ 3)], s08[(d1+ 5)]} <= Sort2(s07[(d1+ 3)], s07[(d1+ 5)]);
        {s08[(d1+ 6)], s08[(d1+ 8)]} <= Sort2(s07[(d1+ 6)], s07[(d1+ 8)]);
        {s08[(d1+ 7)], s08[(d1+ 9)]} <= Sort2(s07[(d1+ 7)], s07[(d1+ 9)]);
        {s08[(d1+10)], s08[(d1+12)]} <= Sort2(s07[(d1+10)], s07[(d1+12)]);
        {s08[(d1+11)], s08[(d1+13)]} <= Sort2(s07[(d1+11)], s07[(d1+13)]);
                    s08[(d1+14)] <= s07[(d1+14)];
                    s08[(d1+15)] <= s07[(d1+15)];

        //stage9
                    s09[(d1+0)] <= s08[(d1+0)];
        {s09[(d1+ 1)], s09[(d1+ 2)]} <= Sort2(s08[(d1+ 1)], s08[(d1+ 2)]);
        {s09[(d1+ 3)], s09[(d1+ 4)]} <= Sort2(s08[(d1+ 3)], s08[(d1+ 4)]);
        {s09[(d1+ 5)], s09[(d1+ 6)]} <= Sort2(s08[(d1+ 5)], s08[(d1+ 6)]);
        {s09[(d1+ 7)], s09[(d1+ 8)]} <= Sort2(s08[(d1+ 7)], s08[(d1+ 8)]);
        {s09[(d1+ 9)], s09[(d1+10)]} <= Sort2(s08[(d1+ 9)], s08[(d1+10)]);
        {s09[(d1+11)], s09[(d1+12)]} <= Sort2(s08[(d1+11)], s08[(d1+12)]);
        {s09[(d1+13)], s09[(d1+14)]} <= Sort2(s08[(d1+13)], s08[(d1+14)]);
                    s09[(d1+15)] <= s08[(d1+15)];
    end
    s06[(48)] <= s05[(48)];
    s07[(48)] <= s06[(48)];
    s08[(48)] <= s07[(48)];
    s09[(48)] <= s08[(48)];

    sr_bypass_data[6] <= sr_bypass_data[5];
    sr_de[6] <= sr_de[5];
    sr_hs[6] <= sr_hs[5];
    sr_vs[6] <= sr_vs[5];

    sr_bypass_data[7] <= sr_bypass_data[6];
    sr_de[7] <= sr_de[6];
    sr_hs[7] <= sr_hs[6];
    sr_vs[7] <= sr_vs[6];

    sr_bypass_data[8] <= sr_bypass_data[7];
    sr_de[8] <= sr_de[7];
    sr_hs[8] <= sr_hs[7];
    sr_vs[8] <= sr_vs[7];

    sr_bypass_data[9] <= sr_bypass_data[8];
    sr_de[9] <= sr_de[8];
    sr_hs[9] <= sr_hs[8];
    sr_vs[9] <= sr_vs[8];

    for (e=0; e<32; e=e+32) begin
        //stage10
        {s10[(e+ 0)], s10[(e+16)]} <= Sort2(s09[(e+ 0)], s09[(e+16)]);
        {s10[(e+ 1)], s10[(e+17)]} <= Sort2(s09[(e+ 1)], s09[(e+17)]);
        {s10[(e+ 2)], s10[(e+18)]} <= Sort2(s09[(e+ 2)], s09[(e+18)]);
        {s10[(e+ 3)], s10[(e+19)]} <= Sort2(s09[(e+ 3)], s09[(e+19)]);
        {s10[(e+ 4)], s10[(e+20)]} <= Sort2(s09[(e+ 4)], s09[(e+20)]);
        {s10[(e+ 5)], s10[(e+21)]} <= Sort2(s09[(e+ 5)], s09[(e+21)]);
        {s10[(e+ 6)], s10[(e+22)]} <= Sort2(s09[(e+ 6)], s09[(e+22)]);
        {s10[(e+ 7)], s10[(e+23)]} <= Sort2(s09[(e+ 7)], s09[(e+23)]);
        {s10[(e+ 8)], s10[(e+24)]} <= Sort2(s09[(e+ 8)], s09[(e+24)]);
        {s10[(e+ 9)], s10[(e+25)]} <= Sort2(s09[(e+ 9)], s09[(e+25)]);
        {s10[(e+10)], s10[(e+26)]} <= Sort2(s09[(e+10)], s09[(e+26)]);
        {s10[(e+11)], s10[(e+27)]} <= Sort2(s09[(e+11)], s09[(e+27)]);
        {s10[(e+12)], s10[(e+28)]} <= Sort2(s09[(e+12)], s09[(e+28)]);
        {s10[(e+13)], s10[(e+29)]} <= Sort2(s09[(e+13)], s09[(e+29)]);
        {s10[(e+14)], s10[(e+30)]} <= Sort2(s09[(e+14)], s09[(e+30)]);
        {s10[(e+15)], s10[(e+31)]} <= Sort2(s09[(e+15)], s09[(e+31)]);

        //stage11
                    s11[(e+0)] <= s10[(e+0)];
                    s11[(e+1)] <= s10[(e+1)];
                    s11[(e+2)] <= s10[(e+2)];
                    s11[(e+3)] <= s10[(e+3)];
                    s11[(e+4)] <= s10[(e+4)];
                    s11[(e+5)] <= s10[(e+5)];
                    s11[(e+6)] <= s10[(e+6)];
                    s11[(e+7)] <= s10[(e+7)];
        {s11[(e+ 8)], s11[(e+16)]} <= Sort2(s10[(e+ 8)], s10[(e+16)]);
        {s11[(e+ 9)], s11[(e+17)]} <= Sort2(s10[(e+ 9)], s10[(e+17)]);
        {s11[(e+10)], s11[(e+18)]} <= Sort2(s10[(e+10)], s10[(e+18)]);
        {s11[(e+11)], s11[(e+19)]} <= Sort2(s10[(e+11)], s10[(e+19)]);
        {s11[(e+12)], s11[(e+20)]} <= Sort2(s10[(e+12)], s10[(e+20)]);
        {s11[(e+13)], s11[(e+21)]} <= Sort2(s10[(e+13)], s10[(e+21)]);
        {s11[(e+14)], s11[(e+22)]} <= Sort2(s10[(e+14)], s10[(e+22)]);
        {s11[(e+15)], s11[(e+23)]} <= Sort2(s10[(e+15)], s10[(e+23)]);
                    s11[(e+24)] <= s10[(e+24)];
                    s11[(e+25)] <= s10[(e+25)];
                    s11[(e+26)] <= s10[(e+26)];
                    s11[(e+27)] <= s10[(e+27)];
                    s11[(e+28)] <= s10[(e+28)];
                    s11[(e+29)] <= s10[(e+29)];
                    s11[(e+30)] <= s10[(e+30)];
                    s11[(e+31)] <= s10[(e+31)];

        //stage12
                    s12[(e+0)] <= s11[(e+0)];
                    s12[(e+1)] <= s11[(e+1)];
                    s12[(e+2)] <= s11[(e+2)];
                    s12[(e+3)] <= s11[(e+3)];
        {s12[(e+ 4)], s12[(e+ 8)]} <= Sort2(s11[(e+ 4)], s11[(e+ 8)]);
        {s12[(e+ 5)], s12[(e+ 9)]} <= Sort2(s11[(e+ 5)], s11[(e+ 9)]);
        {s12[(e+ 6)], s12[(e+10)]} <= Sort2(s11[(e+ 6)], s11[(e+10)]);
        {s12[(e+ 7)], s12[(e+11)]} <= Sort2(s11[(e+ 7)], s11[(e+11)]);
        {s12[(e+12)], s12[(e+16)]} <= Sort2(s11[(e+12)], s11[(e+16)]);
        {s12[(e+13)], s12[(e+17)]} <= Sort2(s11[(e+13)], s11[(e+17)]);
        {s12[(e+14)], s12[(e+18)]} <= Sort2(s11[(e+14)], s11[(e+18)]);
        {s12[(e+15)], s12[(e+19)]} <= Sort2(s11[(e+15)], s11[(e+19)]);
        {s12[(e+20)], s12[(e+24)]} <= Sort2(s11[(e+20)], s11[(e+24)]);
        {s12[(e+21)], s12[(e+25)]} <= Sort2(s11[(e+21)], s11[(e+25)]);
        {s12[(e+22)], s12[(e+26)]} <= Sort2(s11[(e+22)], s11[(e+26)]);
        {s12[(e+23)], s12[(e+27)]} <= Sort2(s11[(e+23)], s11[(e+27)]);
                    s12[(e+28)] <= s11[(e+28)];
                    s12[(e+29)] <= s11[(e+29)];
                    s12[(e+30)] <= s11[(e+30)];
                    s12[(e+31)] <= s11[(e+31)];

        //stage13
                    s13[(e+0)] <= s12[(e+0)];
                    s13[(e+1)] <= s12[(e+1)];
        {s13[(e+ 2)], s13[(e+ 4)]} <= Sort2(s12[(e+ 2)], s12[(e+ 4)]);
        {s13[(e+ 3)], s13[(e+ 5)]} <= Sort2(s12[(e+ 3)], s12[(e+ 5)]);
        {s13[(e+ 6)], s13[(e+ 8)]} <= Sort2(s12[(e+ 6)], s12[(e+ 8)]);
        {s13[(e+ 7)], s13[(e+ 9)]} <= Sort2(s12[(e+ 7)], s12[(e+ 9)]);
        {s13[(e+10)], s13[(e+12)]} <= Sort2(s12[(e+10)], s12[(e+12)]);
        {s13[(e+11)], s13[(e+13)]} <= Sort2(s12[(e+11)], s12[(e+13)]);
        {s13[(e+14)], s13[(e+16)]} <= Sort2(s12[(e+14)], s12[(e+16)]);
        {s13[(e+15)], s13[(e+17)]} <= Sort2(s12[(e+15)], s12[(e+17)]);
        {s13[(e+18)], s13[(e+20)]} <= Sort2(s12[(e+18)], s12[(e+20)]);
        {s13[(e+19)], s13[(e+21)]} <= Sort2(s12[(e+19)], s12[(e+21)]);
        {s13[(e+22)], s13[(e+24)]} <= Sort2(s12[(e+22)], s12[(e+24)]);
        {s13[(e+23)], s13[(e+25)]} <= Sort2(s12[(e+23)], s12[(e+25)]);
        {s13[(e+26)], s13[(e+28)]} <= Sort2(s12[(e+26)], s12[(e+28)]);
        {s13[(e+27)], s13[(e+29)]} <= Sort2(s12[(e+27)], s12[(e+29)]);
                    s13[(e+30)] <= s12[(e+30)];
                    s13[(e+31)] <= s12[(e+31)];

        //stage14
                    s14[(e+0)] <= s13[(e+0)];
        {s14[(e+ 1)], s14[(e+ 2)]} <= Sort2(s13[(e+ 1)], s13[(e+ 2)]);
        {s14[(e+ 3)], s14[(e+ 4)]} <= Sort2(s13[(e+ 3)], s13[(e+ 4)]);
        {s14[(e+ 5)], s14[(e+ 6)]} <= Sort2(s13[(e+ 5)], s13[(e+ 6)]);
        {s14[(e+ 7)], s14[(e+ 8)]} <= Sort2(s13[(e+ 7)], s13[(e+ 8)]);
        {s14[(e+ 9)], s14[(e+10)]} <= Sort2(s13[(e+ 9)], s13[(e+10)]);
        {s14[(e+11)], s14[(e+12)]} <= Sort2(s13[(e+11)], s13[(e+12)]);
        {s14[(e+13)], s14[(e+14)]} <= Sort2(s13[(e+13)], s13[(e+14)]);
        {s14[(e+15)], s14[(e+16)]} <= Sort2(s13[(e+15)], s13[(e+16)]);
        {s14[(e+17)], s14[(e+18)]} <= Sort2(s13[(e+17)], s13[(e+18)]);
        {s14[(e+19)], s14[(e+20)]} <= Sort2(s13[(e+19)], s13[(e+20)]);
        {s14[(e+21)], s14[(e+22)]} <= Sort2(s13[(e+21)], s13[(e+22)]);
        {s14[(e+23)], s14[(e+24)]} <= Sort2(s13[(e+23)], s13[(e+24)]);
        {s14[(e+25)], s14[(e+26)]} <= Sort2(s13[(e+25)], s13[(e+26)]);
        {s14[(e+27)], s14[(e+28)]} <= Sort2(s13[(e+27)], s13[(e+28)]);
        {s14[(e+29)], s14[(e+30)]} <= Sort2(s13[(e+29)], s13[(e+30)]);
                    s14[(e+31)] <= s13[(e+31)];
    end
    //stage10
    {s10[(32)], s10[(48)]} <= Sort2(s09[(32)], s09[(48)]);
    s10[(33)] <= s09[(33)];
    s10[(34)] <= s09[(34)];
    s10[(35)] <= s09[(35)];
    s10[(36)] <= s09[(36)];
    s10[(37)] <= s09[(37)];
    s10[(38)] <= s09[(38)];
    s10[(39)] <= s09[(39)];
    s10[(40)] <= s09[(40)];
    s10[(41)] <= s09[(41)];
    s10[(42)] <= s09[(42)];
    s10[(43)] <= s09[(43)];
    s10[(44)] <= s09[(44)];
    s10[(45)] <= s09[(45)];
    s10[(46)] <= s09[(46)];
    s10[(47)] <= s09[(47)];

    sr_bypass_data[10] <= sr_bypass_data[9];
    sr_de[10] <= sr_de[9];
    sr_hs[10] <= sr_hs[9];
    sr_vs[10] <= sr_vs[9];

    //stage11
    s11[(32)] <= s10[(32)];
    s11[(33)] <= s10[(33)];
    s11[(34)] <= s10[(34)];
    s11[(35)] <= s10[(35)];
    s11[(36)] <= s10[(36)];
    s11[(37)] <= s10[(37)];
    s11[(38)] <= s10[(38)];
    s11[(39)] <= s10[(39)];
    {s11[(40)], s11[(48)]} <= Sort2(s10[(40)], s10[(48)]);
    s11[(41)] <= s10[(41)];
    s11[(42)] <= s10[(42)];
    s11[(43)] <= s10[(43)];
    s11[(44)] <= s10[(44)];
    s11[(45)] <= s10[(45)];
    s11[(46)] <= s10[(46)];
    s11[(47)] <= s10[(47)];

    sr_bypass_data[11] <= sr_bypass_data[10];
    sr_de[11] <= sr_de[10];
    sr_hs[11] <= sr_hs[10];
    sr_vs[11] <= sr_vs[10];

    //stage12
    s12[(32)] <= s11[(32)];
    s12[(33)] <= s11[(33)];
    s12[(34)] <= s11[(34)];
    s12[(35)] <= s11[(35)];
    {s12[(36)], s12[(40)]} <= Sort2(s11[(36)], s11[(40)]);
    {s12[(37)], s12[(41)]} <= Sort2(s11[(37)], s11[(41)]);
    {s12[(38)], s12[(42)]} <= Sort2(s11[(38)], s11[(42)]);
    {s12[(39)], s12[(43)]} <= Sort2(s11[(39)], s11[(43)]);
    {s12[(44)], s12[(48)]} <= Sort2(s11[(44)], s11[(48)]);
    s12[(45)] <= s11[(45)];
    s12[(46)] <= s11[(46)];
    s12[(47)] <= s11[(47)];

    sr_bypass_data[12] <= sr_bypass_data[11];
    sr_de[12] <= sr_de[11];
    sr_hs[12] <= sr_hs[11];
    sr_vs[12] <= sr_vs[11];

    //stage13
    s13[(32)] <= s12[(32)];
    s13[(33)] <= s12[(33)];
    {s13[(34)], s13[(36)]} <= Sort2(s12[(34)], s12[(36)]);
    {s13[(35)], s13[(37)]} <= Sort2(s12[(35)], s12[(37)]);
    {s13[(38)], s13[(40)]} <= Sort2(s12[(38)], s12[(40)]);
    {s13[(39)], s13[(41)]} <= Sort2(s12[(39)], s12[(41)]);
    {s13[(42)], s13[(44)]} <= Sort2(s12[(42)], s12[(44)]);
    {s13[(43)], s13[(45)]} <= Sort2(s12[(43)], s12[(45)]);
    {s13[(46)], s13[(48)]} <= Sort2(s12[(46)], s12[(48)]);
    s13[(47)] <= s12[(47)];

    sr_bypass_data[13] <= sr_bypass_data[12];
    sr_de[13] <= sr_de[12];
    sr_hs[13] <= sr_hs[12];
    sr_vs[13] <= sr_vs[12];

    //stage14
    s14[(32)] <= s13[(32)];
    {s14[(33)], s14[(34)]} <= Sort2(s13[(33)], s13[(34)]);
    {s14[(35)], s14[(36)]} <= Sort2(s13[(35)], s13[(36)]);
    {s14[(37)], s14[(38)]} <= Sort2(s13[(37)], s13[(38)]);
    {s14[(39)], s14[(40)]} <= Sort2(s13[(39)], s13[(40)]);
    {s14[(41)], s14[(42)]} <= Sort2(s13[(41)], s13[(42)]);
    {s14[(43)], s14[(44)]} <= Sort2(s13[(43)], s13[(44)]);
    {s14[(45)], s14[(46)]} <= Sort2(s13[(45)], s13[(46)]);
    {s14[(47)], s14[(48)]} <= Sort2(s13[(47)], s13[(48)]);

    sr_bypass_data[14] <= sr_bypass_data[13];
    sr_de[14] <= sr_de[13];
    sr_hs[14] <= sr_hs[13];
    sr_vs[14] <= sr_vs[13];

    //stage15
    {s15[( 0)], s15[(32)]} <= Sort2(s14[( 0)], s14[(32)]);
    {s15[( 1)], s15[(33)]} <= Sort2(s14[( 1)], s14[(33)]);
    {s15[( 2)], s15[(34)]} <= Sort2(s14[( 2)], s14[(34)]);
    {s15[( 3)], s15[(35)]} <= Sort2(s14[( 3)], s14[(35)]);
    {s15[( 4)], s15[(36)]} <= Sort2(s14[( 4)], s14[(36)]);
    {s15[( 5)], s15[(37)]} <= Sort2(s14[( 5)], s14[(37)]);
    {s15[( 6)], s15[(38)]} <= Sort2(s14[( 6)], s14[(38)]);
    {s15[( 7)], s15[(39)]} <= Sort2(s14[( 7)], s14[(39)]);
    {s15[( 8)], s15[(40)]} <= Sort2(s14[( 8)], s14[(40)]);
    {s15[( 9)], s15[(41)]} <= Sort2(s14[( 9)], s14[(41)]);
    {s15[(10)], s15[(42)]} <= Sort2(s14[(10)], s14[(42)]);
    {s15[(11)], s15[(43)]} <= Sort2(s14[(11)], s14[(43)]);
    {s15[(12)], s15[(44)]} <= Sort2(s14[(12)], s14[(44)]);
    {s15[(13)], s15[(45)]} <= Sort2(s14[(13)], s14[(45)]);
    {s15[(14)], s15[(46)]} <= Sort2(s14[(14)], s14[(46)]);
    {s15[(15)], s15[(47)]} <= Sort2(s14[(15)], s14[(47)]);
    {s15[(16)], s15[(48)]} <= Sort2(s14[(16)], s14[(48)]);
    s15[(17)] <= s14[(17)];
    s15[(18)] <= s14[(18)];
    s15[(19)] <= s14[(19)];
    s15[(20)] <= s14[(20)];
    s15[(21)] <= s14[(21)];
    s15[(22)] <= s14[(22)];
    s15[(23)] <= s14[(23)];
    s15[(24)] <= s14[(24)];
    s15[(25)] <= s14[(25)];
    s15[(26)] <= s14[(26)];
    s15[(27)] <= s14[(27)];
    s15[(28)] <= s14[(28)];
    s15[(29)] <= s14[(29)];
    s15[(30)] <= s14[(30)];
    s15[(31)] <= s14[(31)];

    sr_bypass_data[15] <= sr_bypass_data[14];
    sr_de[15] <= sr_de[14];
    sr_hs[15] <= sr_hs[14];
    sr_vs[15] <= sr_vs[14];

    //stage16
    s16[( 0)] <= s15[( 0)];
    s16[( 1)] <= s15[( 1)];
    s16[( 2)] <= s15[( 2)];
    s16[( 3)] <= s15[( 3)];
    s16[( 4)] <= s15[( 4)];
    s16[( 5)] <= s15[( 5)];
    s16[( 6)] <= s15[( 6)];
    s16[( 7)] <= s15[( 7)];
    s16[( 8)] <= s15[( 8)];
    s16[( 9)] <= s15[( 9)];
    s16[(10)] <= s15[(10)];
    s16[(11)] <= s15[(11)];
    s16[(12)] <= s15[(12)];
    s16[(13)] <= s15[(13)];
    s16[(14)] <= s15[(14)];
    s16[(15)] <= s15[(15)];
    {s16[(16)], s16[(32)]} <= Sort2(s15[(16)], s15[(32)]);
    {s16[(17)], s16[(33)]} <= Sort2(s15[(17)], s15[(33)]);
    {s16[(18)], s16[(34)]} <= Sort2(s15[(18)], s15[(34)]);
    {s16[(19)], s16[(35)]} <= Sort2(s15[(19)], s15[(35)]);
    {s16[(20)], s16[(36)]} <= Sort2(s15[(20)], s15[(36)]);
    {s16[(21)], s16[(37)]} <= Sort2(s15[(21)], s15[(37)]);
    {s16[(22)], s16[(38)]} <= Sort2(s15[(22)], s15[(38)]);
    {s16[(23)], s16[(39)]} <= Sort2(s15[(23)], s15[(39)]);
    {s16[(24)], s16[(40)]} <= Sort2(s15[(24)], s15[(40)]);
    {s16[(25)], s16[(41)]} <= Sort2(s15[(25)], s15[(41)]);
    {s16[(26)], s16[(42)]} <= Sort2(s15[(26)], s15[(42)]);
    {s16[(27)], s16[(43)]} <= Sort2(s15[(27)], s15[(43)]);
    {s16[(28)], s16[(44)]} <= Sort2(s15[(28)], s15[(44)]);
    {s16[(29)], s16[(45)]} <= Sort2(s15[(29)], s15[(45)]);
    {s16[(30)], s16[(46)]} <= Sort2(s15[(30)], s15[(46)]);
    {s16[(31)], s16[(47)]} <= Sort2(s15[(31)], s15[(47)]);
    s16[(48)] <= s15[(48)];

    sr_bypass_data[16] <= sr_bypass_data[15];
    sr_de[16] <= sr_de[15];
    sr_hs[16] <= sr_hs[15];
    sr_vs[16] <= sr_vs[15];

    //stage17
    s17[(0)] <= s16[(0)];
    s17[(1)] <= s16[(1)];
    s17[(2)] <= s16[(2)];
    s17[(3)] <= s16[(3)];
    s17[(4)] <= s16[(4)];
    s17[(5)] <= s16[(5)];
    s17[(6)] <= s16[(6)];
    s17[(7)] <= s16[(7)];

    {s17[( 8)], s17[(16)]} <= Sort2(s16[( 8)], s16[(16)]);
    {s17[( 9)], s17[(17)]} <= Sort2(s16[( 9)], s16[(17)]);
    {s17[(10)], s17[(18)]} <= Sort2(s16[(10)], s16[(18)]);
    {s17[(11)], s17[(19)]} <= Sort2(s16[(11)], s16[(19)]);
    {s17[(12)], s17[(20)]} <= Sort2(s16[(12)], s16[(20)]);
    {s17[(13)], s17[(21)]} <= Sort2(s16[(13)], s16[(21)]);
    {s17[(14)], s17[(22)]} <= Sort2(s16[(14)], s16[(22)]);
    {s17[(15)], s17[(23)]} <= Sort2(s16[(15)], s16[(23)]);

    {s17[(24)], s17[(32)]} <= Sort2(s16[(24)], s16[(32)]);
    {s17[(25)], s17[(33)]} <= Sort2(s16[(25)], s16[(33)]);
    {s17[(26)], s17[(34)]} <= Sort2(s16[(26)], s16[(34)]);
    {s17[(27)], s17[(35)]} <= Sort2(s16[(27)], s16[(35)]);
    {s17[(28)], s17[(36)]} <= Sort2(s16[(28)], s16[(36)]);
    {s17[(29)], s17[(37)]} <= Sort2(s16[(29)], s16[(37)]);
    {s17[(30)], s17[(38)]} <= Sort2(s16[(30)], s16[(38)]);
    {s17[(31)], s17[(39)]} <= Sort2(s16[(31)], s16[(39)]);

    {s17[(40)], s17[(48)]} <= Sort2(s16[(40)], s16[(48)]);

    s17[(41)] <= s16[(41)];
    s17[(42)] <= s16[(42)];
    s17[(43)] <= s16[(43)];
    s17[(44)] <= s16[(44)];
    s17[(45)] <= s16[(45)];
    s17[(46)] <= s16[(46)];
    s17[(47)] <= s16[(47)];

    sr_bypass_data[17] <= sr_bypass_data[16];
    sr_de[17] <= sr_de[16];
    sr_hs[17] <= sr_hs[16];
    sr_vs[17] <= sr_vs[16];

    //stage18
    s18[(0)] <= s17[(0)];
    s18[(1)] <= s17[(1)];
    s18[(2)] <= s17[(2)];
    s18[(3)] <= s17[(3)];

    {s18[( 4)], s18[( 8)]} <= Sort2(s17[( 4)], s17[( 8)]);
    {s18[( 5)], s18[( 9)]} <= Sort2(s17[( 5)], s17[( 9)]);
    {s18[( 6)], s18[(10)]} <= Sort2(s17[( 6)], s17[(10)]);
    {s18[( 7)], s18[(11)]} <= Sort2(s17[( 7)], s17[(11)]);

    {s18[(12)], s18[(16)]} <= Sort2(s17[(12)], s17[(16)]);
    {s18[(13)], s18[(17)]} <= Sort2(s17[(13)], s17[(17)]);
    {s18[(14)], s18[(18)]} <= Sort2(s17[(14)], s17[(18)]);
    {s18[(15)], s18[(19)]} <= Sort2(s17[(15)], s17[(19)]);

    {s18[(20)], s18[(24)]} <= Sort2(s17[(20)], s17[(24)]);
    {s18[(21)], s18[(25)]} <= Sort2(s17[(21)], s17[(25)]);
    {s18[(22)], s18[(26)]} <= Sort2(s17[(22)], s17[(26)]);
    {s18[(23)], s18[(27)]} <= Sort2(s17[(23)], s17[(27)]);

    {s18[(28)], s18[(32)]} <= Sort2(s17[(28)], s17[(32)]);
    {s18[(29)], s18[(33)]} <= Sort2(s17[(29)], s17[(33)]);
    {s18[(30)], s18[(34)]} <= Sort2(s17[(30)], s17[(34)]);
    {s18[(31)], s18[(35)]} <= Sort2(s17[(31)], s17[(35)]);

    {s18[(36)], s18[(40)]} <= Sort2(s17[(36)], s17[(40)]);
    {s18[(37)], s18[(41)]} <= Sort2(s17[(37)], s17[(41)]);
    {s18[(38)], s18[(42)]} <= Sort2(s17[(38)], s17[(42)]);
    {s18[(39)], s18[(43)]} <= Sort2(s17[(39)], s17[(43)]);

    {s18[(44)], s18[(48)]} <= Sort2(s17[(44)], s17[(48)]);

    s18[(45)] <= s17[(45)];
    s18[(46)] <= s17[(46)];
    s18[(47)] <= s17[(47)];

    sr_bypass_data[18] <= sr_bypass_data[17];
    sr_de[18] <= sr_de[17];
    sr_hs[18] <= sr_hs[17];
    sr_vs[18] <= sr_vs[17];

    //stage19
    s19[(0)] <= s18[(0)];
    s19[(1)] <= s18[(1)];

    {s19[( 2)], s19[( 4)]} <= Sort2(s18[( 2)], s18[( 4)]);
    {s19[( 3)], s19[( 5)]} <= Sort2(s18[( 3)], s18[( 5)]);

    {s19[( 6)], s19[( 8)]} <= Sort2(s18[( 6)], s18[( 8)]);
    {s19[( 7)], s19[( 9)]} <= Sort2(s18[( 7)], s18[( 9)]);

    {s19[(10)], s19[(12)]} <= Sort2(s18[(10)], s18[(12)]);
    {s19[(11)], s19[(13)]} <= Sort2(s18[(11)], s18[(13)]);

    {s19[(14)], s19[(16)]} <= Sort2(s18[(14)], s18[(16)]);
    {s19[(15)], s19[(17)]} <= Sort2(s18[(15)], s18[(17)]);

    {s19[(18)], s19[(20)]} <= Sort2(s18[(18)], s18[(20)]);
    {s19[(19)], s19[(21)]} <= Sort2(s18[(19)], s18[(21)]);

    {s19[(22)], s19[(24)]} <= Sort2(s18[(22)], s18[(24)]);
    {s19[(23)], s19[(25)]} <= Sort2(s18[(23)], s18[(25)]);

    {s19[(26)], s19[(28)]} <= Sort2(s18[(26)], s18[(28)]);
    {s19[(27)], s19[(29)]} <= Sort2(s18[(27)], s18[(29)]);

    {s19[(30)], s19[(32)]} <= Sort2(s18[(30)], s18[(32)]);
    {s19[(31)], s19[(33)]} <= Sort2(s18[(31)], s18[(33)]);

    {s19[(34)], s19[(36)]} <= Sort2(s18[(34)], s18[(36)]);
    {s19[(35)], s19[(37)]} <= Sort2(s18[(35)], s18[(37)]);

    {s19[(38)], s19[(40)]} <= Sort2(s18[(38)], s18[(40)]);
    {s19[(39)], s19[(41)]} <= Sort2(s18[(39)], s18[(41)]);

    {s19[(42)], s19[(44)]} <= Sort2(s18[(42)], s18[(44)]);
    {s19[(43)], s19[(45)]} <= Sort2(s18[(43)], s18[(45)]);

    {s19[(46)], s19[(48)]} <= Sort2(s18[(46)], s18[(48)]);
    s19[(47)] <= s18[(47)];

    sr_bypass_data[19] <= sr_bypass_data[18];
    sr_de[19] <= sr_de[18];
    sr_hs[19] <= sr_hs[18];
    sr_vs[19] <= sr_vs[18];

    //stage20
    s20[(0)] <= s19[(0)];
    {s20[( 1)], s20[( 2)]} <= Sort2(s19[( 1)], s19[( 2)]);
    {s20[( 3)], s20[( 4)]} <= Sort2(s19[( 3)], s19[( 4)]);
    {s20[( 5)], s20[( 6)]} <= Sort2(s19[( 5)], s19[( 6)]);
    {s20[( 7)], s20[( 8)]} <= Sort2(s19[( 7)], s19[( 8)]);
    {s20[( 9)], s20[(10)]} <= Sort2(s19[( 9)], s19[(10)]);
    {s20[(11)], s20[(12)]} <= Sort2(s19[(11)], s19[(12)]);
    {s20[(13)], s20[(14)]} <= Sort2(s19[(13)], s19[(14)]);
    {s20[(15)], s20[(16)]} <= Sort2(s19[(15)], s19[(16)]);
    {s20[(17)], s20[(18)]} <= Sort2(s19[(17)], s19[(18)]);
    {s20[(19)], s20[(20)]} <= Sort2(s19[(19)], s19[(20)]);
    {s20[(21)], s20[(22)]} <= Sort2(s19[(21)], s19[(22)]);
    {s20[(23)], s20[(24)]} <= Sort2(s19[(23)], s19[(24)]);
    {s20[(25)], s20[(26)]} <= Sort2(s19[(25)], s19[(26)]);
    {s20[(27)], s20[(28)]} <= Sort2(s19[(27)], s19[(28)]);
    {s20[(29)], s20[(30)]} <= Sort2(s19[(29)], s19[(30)]);
    {s20[(31)], s20[(32)]} <= Sort2(s19[(31)], s19[(32)]);
    {s20[(33)], s20[(34)]} <= Sort2(s19[(33)], s19[(34)]);
    {s20[(35)], s20[(36)]} <= Sort2(s19[(35)], s19[(36)]);
    {s20[(37)], s20[(38)]} <= Sort2(s19[(37)], s19[(38)]);
    {s20[(39)], s20[(40)]} <= Sort2(s19[(39)], s19[(40)]);
    {s20[(41)], s20[(42)]} <= Sort2(s19[(41)], s19[(42)]);
    {s20[(43)], s20[(44)]} <= Sort2(s19[(43)], s19[(44)]);
    {s20[(45)], s20[(46)]} <= Sort2(s19[(45)], s19[(46)]);
    {s20[(47)], s20[(48)]} <= Sort2(s19[(47)], s19[(48)]);

    sr_bypass_data[20] <= sr_bypass_data[19];
    sr_de[20] <= sr_de[19];
    sr_hs[20] <= sr_hs[19];
    sr_vs[20] <= sr_vs[19];
end

genvar k;
generate
    for (k=0; k<KERNEL_SIZE; k=k+1) begin
        assign xo[k*8 +: PIXEL_WIDTH] = s20[k];
    end
endgenerate

assign do_o = s20[(24)];
assign de_o = sr_de[20];
assign hs_o = sr_hs[20];
assign vs_o = sr_vs[20];
assign bypass_o = sr_bypass_data[20];

endmodule


