-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor + Kukla Anatol
--
-- Create Date : 18.01.2012 17:24:28
-- Module Name : hdd_main
--
-- ����������/�������� :
--
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.vicg_common_pkg.all;
use work.prj_cfg.all;
use work.cfgdev_pkg.all;
use work.sata_glob_pkg.all;
use work.dsn_hdd_pkg.all;
use work.hdd_main_unit_pkg.all;
use work.video_ctrl_pkg.all;
use work.mem_ctrl_pkg.all;

entity hdd_main is
generic(
G_VSYN_ACTIVE : std_logic:='1';
G_SIM : string:="OFF"
);
port(
--------------------------------------------------
--VideoIN
--------------------------------------------------
p_in_vd       : in   std_logic_vector(99 downto 0);
p_in_vin_vs   : in   std_logic;
p_in_vin_hs   : in   std_logic;
p_in_vin_clk  : in   std_logic;

--------------------------------------------------
--VideoOUT
--------------------------------------------------
p_out_vd      : out  std_logic_vector(31 downto 0);
p_in_vout_vs  : in   std_logic;
p_in_vout_hs  : in   std_logic;
p_in_vout_clk : in   std_logic;

--------------------------------------------------
--RAM
--------------------------------------------------
p_out_mcb5_a        : out   std_logic_vector(12 downto 0);--(C5_MEM_ADDR_WIDTH-1 downto 0);
p_out_mcb5_ba       : out   std_logic_vector(2 downto 0) ;--(C5_MEM_BANKADDR_WIDTH-1 downto 0);
p_out_mcb5_ras_n    : out   std_logic;
p_out_mcb5_cas_n    : out   std_logic;
p_out_mcb5_we_n     : out   std_logic;
p_out_mcb5_odt      : out   std_logic;
p_out_mcb5_cke      : out   std_logic;
p_out_mcb5_dm       : out   std_logic;
p_out_mcb5_udm      : out   std_logic;
p_out_mcb5_ck       : out   std_logic;
p_out_mcb5_ck_n     : out   std_logic;
p_inout_mcb5_dq     : inout std_logic_vector(15 downto 0);--(C5_NUM_DQ_PINS-1 downto 0);
p_inout_mcb5_udqs   : inout std_logic;
p_inout_mcb5_udqs_n : inout std_logic;
p_inout_mcb5_dqs    : inout std_logic;
p_inout_mcb5_dqs_n  : inout std_logic;
p_inout_mcb5_rzq    : inout std_logic;
p_inout_mcb5_zio    : inout std_logic;

p_out_mcb1_a        : out   std_logic_vector(12 downto 0);--(C5_MEM_ADDR_WIDTH-1 downto 0);
p_out_mcb1_ba       : out   std_logic_vector(2 downto 0) ;--(C5_MEM_BANKADDR_WIDTH-1 downto 0);
p_out_mcb1_ras_n    : out   std_logic;
p_out_mcb1_cas_n    : out   std_logic;
p_out_mcb1_we_n     : out   std_logic;
p_out_mcb1_odt      : out   std_logic;
p_out_mcb1_cke      : out   std_logic;
p_out_mcb1_dm       : out   std_logic;
p_out_mcb1_udm      : out   std_logic;
p_out_mcb1_ck       : out   std_logic;
p_out_mcb1_ck_n     : out   std_logic;
p_inout_mcb1_dq     : inout std_logic_vector(15 downto 0);--(C5_NUM_DQ_PINS-1 downto 0);
p_inout_mcb1_udqs   : inout std_logic;
p_inout_mcb1_udqs_n : inout std_logic;
p_inout_mcb1_dqs    : inout std_logic;
p_inout_mcb1_dqs_n  : inout std_logic;
p_inout_mcb1_rzq    : inout std_logic;
p_inout_mcb1_zio    : inout std_logic;

--------------------------------------------------
--SATA
--------------------------------------------------
p_out_sata_txn      : out   std_logic_vector((C_SH_GTCH_COUNT_MAX*C_SH_COUNT_MAX(C_PCFG_HDD_COUNT-1))-1 downto 0);--std_logic_vector(3 downto 0);
p_out_sata_txp      : out   std_logic_vector((C_SH_GTCH_COUNT_MAX*C_SH_COUNT_MAX(C_PCFG_HDD_COUNT-1))-1 downto 0);--std_logic_vector(3 downto 0);
p_in_sata_rxn       : in    std_logic_vector((C_SH_GTCH_COUNT_MAX*C_SH_COUNT_MAX(C_PCFG_HDD_COUNT-1))-1 downto 0);--std_logic_vector(3 downto 0);
p_in_sata_rxp       : in    std_logic_vector((C_SH_GTCH_COUNT_MAX*C_SH_COUNT_MAX(C_PCFG_HDD_COUNT-1))-1 downto 0);--std_logic_vector(3 downto 0);
p_in_sata_clk_n     : in    std_logic_vector(0 downto 0);
p_in_sata_clk_p     : in    std_logic_vector(0 downto 0);

--------------------------------------------------
--System
--------------------------------------------------
p_out_hdd_grefclk150M : out   std_logic;

p_out_hdd_dcm_lock    : out   std_logic;
p_out_hdd_dcm_gclk75M : out   std_logic;
p_out_hdd_dcm_gclk300M: out   std_logic;
p_out_hdd_dcm_gclk150M: out   std_logic;

p_out_hdd_mem_plllock : out   std_logic;
p_out_hdd_mem_gclk375M: out   std_logic;

--------------------------------------------------
--��������������� ����
--------------------------------------------------
p_inout_ftdi_d   : inout std_logic_vector(7 downto 0);
p_out_ftdi_rd_n  : out   std_logic;
p_out_ftdi_wr_n  : out   std_logic;
p_in_ftdi_txe_n  : in    std_logic;
p_in_ftdi_rxf_n  : in    std_logic;
p_in_ftdi_pwren_n: in    std_logic;

p_out_TP         : out   std_logic_vector(7 downto 0);
p_out_led        : out   std_logic_vector(7 downto 0)
);
end entity;

architecture struct of hdd_main is

component dbgcs_iconx1
  PORT (
    CONTROL0 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0));
--    CONTROL1 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0));

end component;

component dbgcs_iconx2
  PORT (
    CONTROL0 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CONTROL1 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0));

end component;

component dbgcs_iconx3
  PORT (
    CONTROL0 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CONTROL1 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CONTROL2 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0));

end component;

component dbgcs_sata_layer
  PORT (
    CONTROL : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CLK : IN STD_LOGIC;
    DATA : IN STD_LOGIC_VECTOR(122 DOWNTO 0);
    TRIG0 : IN STD_LOGIC_VECTOR(41 DOWNTO 0)
    );
end component;

component dbgcs_sata_raid
  PORT (
    CONTROL : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CLK : IN STD_LOGIC;
    DATA : IN STD_LOGIC_VECTOR(172 downto 0); --(122 DOWNTO 0);
    TRIG0 : IN STD_LOGIC_VECTOR(41 DOWNTO 0)
    );
end component;

signal i_dbgcs_sh0_spd                  : std_logic_vector(35 downto 0);
signal i_dbgcs_hdd0_layer               : std_logic_vector(35 downto 0);
signal i_dbgcs_hdd1_layer               : std_logic_vector(35 downto 0);
signal i_dbgcs_hdd_raid                 : std_logic_vector(35 downto 0);
signal i_dbgcs_cfg                      : std_logic_vector(35 downto 0);

signal i_hdd0layer_dbgcs                : TSH_ila;
signal i_hdd1layer_dbgcs                : TSH_ila;
signal i_cfg_dbgcs                      : TSH_ila;
signal i_hddraid_dbgcs                  : TSH_ila;

component hdd_ram_hfifo
port(
din         : in std_logic_vector(31 downto 0);
wr_en       : in std_logic;
wr_clk      : in std_logic;

dout        : out std_logic_vector(31 downto 0);
rd_en       : in std_logic;
rd_clk      : in std_logic;

full        : out std_logic;
almost_full : out std_logic;
empty       : out std_logic;

--clk         : in std_logic;
rst         : in std_logic
);
end component;

constant CI_MEM_AWIDTH : integer:=32;
constant CI_MEM_DWIDTH : integer:=32;

signal i_vfr_prm                        : TFrXY;

signal i_vbufin_dout                    : std_logic_vector(31 downto 0);
signal i_vbufin_rd                      : std_logic;
signal i_vbufin_empty                   : std_logic;
signal i_vbufout_din                    : std_logic_vector(31 downto 0);
signal i_vbufout_wr                     : std_logic;
signal i_vbufout_full                   : std_logic;

signal i_mem_ctrl_rst                   : std_logic;
signal i_mem_ctrl_rdy                   : std_logic_vector(C_MEM_BANK_COUNT-1 downto 0);
signal i_memch0_in_bank                 : TMemINBank;
signal i_memch0_out_bank                : TMemOUTBank;
signal i_memch1_in_bank                 : TMemINBank;
signal i_memch1_out_bank                : TMemOUTBank;

signal i_phymem_out                     : TRam_outs;
signal i_phymem_inout                   : TRam_inouts;

signal i_usrpll_rst                     : std_logic;
signal i_usrpll_lock                    : std_logic;
signal g_memclk                         : std_logic;

signal i_vctrl_rst                      : std_logic;
signal i_sys_rst_cnt                    : std_logic_vector(5 downto 0):=(others=>'0');
signal i_sys_rst                        : std_logic:='0';
signal g_sata_refclkout                 : std_logic;

signal i_hdd_rst                        : std_logic;
signal i_hdd_gt_refclk150               : std_logic_vector(C_SH_COUNT_MAX(C_PCFG_HDD_COUNT-1)-1 downto 0);
signal g_hdd_gt_refclkout               : std_logic;
signal i_hdd_gt_plldet                  : std_logic;
signal i_hdd_dcm_lock                   : std_logic;
signal g_hdd_dcm_gclk75M                : std_logic;--p_out_hdd_dcm_gclk75M,--i_hdd_dcm_gclk2div,
signal g_hdd_dcm_gclk300M               : std_logic;--p_out_hdd_dcm_gclk300M,--i_hdd_dcm_gclk2x,
signal g_hdd_dcm_gclk150M               : std_logic;--p_out_hdd_dcm_gclk300M,--i_hdd_dcm_gclk2x,

signal i_hdd_rbuf_cfg                   : THDDRBufCfg;
signal i_hdd_rbuf_status                : THDDRBufStatus;

signal i_hdd_txdata                     : std_logic_vector(31 downto 0);
signal i_hdd_txdata_wd                  : std_logic;
signal i_hdd_txbuf_full                 : std_logic;
signal i_hdd_txbuf_pfull                : std_logic;
signal i_hdd_txbuf_empty                : std_logic;

signal i_hdd_rxdata                     : std_logic_vector(31 downto 0);
signal i_hdd_rxdata_rd                  : std_logic;
signal i_hdd_rxbuf_empty                : std_logic;
signal i_hdd_rxbuf_pempty               : std_logic;

signal i_dev_adr                        : std_logic_vector(C_CFGPKT_DADR_M_BIT-C_CFGPKT_DADR_L_BIT downto 0);
signal i_cfg_adr                        : std_logic_vector(C_CFGPKT_RADR_M_BIT-C_CFGPKT_RADR_L_BIT downto 0);
signal i_cfg_adr_ld                     : std_logic;
signal i_cfg_adr_fifo                   : std_logic;
signal i_cfg_wd                         : std_logic;
signal i_cfg_rd                         : std_logic;
signal i_cfg_txd                        : std_logic_vector(15 downto 0);
signal i_cfg_rxd                        : std_logic_vector(15 downto 0);
signal i_cfg_txrdy                      : std_logic;
signal i_cfg_rxrdy                      : std_logic;
signal i_cfg_done                       : std_logic;
--signal i_cfg_tstout                     : std_logic_vector(31 downto 0);

signal i_hdd_module_rdy                 : std_logic;
signal i_hdd_module_error               : std_logic;
signal i_hdd_busy                       : std_logic;
--signal i_hdd_hirq                       : std_logic;
signal i_hdd_done                       : std_logic;

signal i_hdd_dbgcs                      : TSH_dbgcs_exp;
signal i_hdd_dbgled                     : THDDLed_SHCountMax;

--signal i_hdd_sim_gt_txdata              : TBus32_SHCountMax;
--signal i_hdd_sim_gt_txcharisk           : TBus04_SHCountMax;
--signal i_hdd_sim_gt_txcomstart          : std_logic_vector(C_HDD_COUNT_MAX-1 downto 0);
signal i_hdd_sim_gt_rxdata              : TBus32_SHCountMax;
signal i_hdd_sim_gt_rxcharisk           : TBus04_SHCountMax;
signal i_hdd_sim_gt_rxstatus            : TBus03_SHCountMax;
signal i_hdd_sim_gt_rxelecidle          : std_logic_vector(C_HDD_COUNT_MAX-1 downto 0);
signal i_hdd_sim_gt_rxdisperr           : TBus04_SHCountMax;
signal i_hdd_sim_gt_rxnotintable        : TBus04_SHCountMax;
signal i_hdd_sim_gt_rxbyteisaligned     : std_logic_vector(C_HDD_COUNT_MAX-1 downto 0);
--signal i_hdd_sim_gt_sim_rst             : std_logic_vector(C_HDD_COUNT_MAX-1 downto 0);
--signal i_hdd_sim_gt_sim_clk             : std_logic_vector(C_HDD_COUNT_MAX-1 downto 0);
--signal i_hdd_tst_in                     : std_logic_vector(31 downto 0);
signal i_hdd_tst_out                    : std_logic_vector(31 downto 0);

signal i_ram_txbuf_full                 : std_logic;
signal i_ram_txbuf_afull                : std_logic;
signal i_ram_txbuf_empty                : std_logic;
signal i_ram_rxbuf_full                 : std_logic;
signal i_ram_rxbuf_afull                : std_logic;
signal i_ram_rxbuf_empty                : std_logic;
signal i_ram_reset_buf                  : std_logic;

signal i_ram_txbuf_rd                   : std_logic;
signal i_ram_rxbuf_wr                   : std_logic;
signal i_ram_rxbuf_din                  : std_logic_vector(31 downto 0);

signal i_test01_led                     : std_logic;
signal i_test02_led                     : std_logic;

signal tst_vctrl_out                    : std_logic_vector(31 downto 0);
signal sr_vctrl_rst                     : std_logic_vector(1 downto 0):=(others=>'0');
signal tst_syn                          : std_logic:='0';

signal i_vin_dout                       : std_logic_vector(31 downto 0);
signal tst_vin_vs                       : std_logic;
signal tst_vin_hs                       : std_logic;
signal tst_vout_vs                      : std_logic;
signal tst_vout_hs                      : std_logic;

signal t_vbufin_rd                      : std_logic;
signal t_vbufin_empty                   : std_logic;



--//MAIN
begin


--***********************************************************
--
--***********************************************************
p_out_hdd_grefclk150M<=g_sata_refclkout;

p_out_hdd_dcm_lock    <=i_hdd_dcm_lock;
p_out_hdd_dcm_gclk75M <=g_hdd_dcm_gclk75M;
p_out_hdd_dcm_gclk300M<=g_hdd_dcm_gclk300M;
p_out_hdd_dcm_gclk150M<=g_hdd_dcm_gclk150M;

p_out_hdd_mem_plllock <='0';--i_usrpll_lock;
p_out_hdd_mem_gclk375M<='0';--g_memclk;


g_memclk<=g_hdd_dcm_gclk300M;
--g_sata_refclkout<=p_in_sata_clk_p(0);

--***********************************************************
--RESET
--***********************************************************
process(g_sata_refclkout)
begin
  if g_sata_refclkout'event and g_sata_refclkout = '1' then
    if i_sys_rst_cnt(i_sys_rst_cnt'high) = '0' then
      i_sys_rst_cnt <= i_sys_rst_cnt + 1;
    end if;
  end if;
end process;

i_sys_rst <= i_sys_rst_cnt(i_sys_rst_cnt'high - 1);
i_hdd_rst <= i_sys_rst;-- or i_hdd_rbuf_cfg.greset;
i_ram_reset_buf<=i_hdd_rst or i_hdd_rbuf_cfg.dmacfg.clr_err;
i_vctrl_rst<= i_sys_rst or not (AND_reduce(i_mem_ctrl_rdy));
i_mem_ctrl_rst <= not i_hdd_dcm_lock or i_hdd_rbuf_cfg.greset;--i_usrpll_lock;--


--***********************************************************
--VIDEO IN/OUT
--***********************************************************
--Video Input
m_vin_cam : vin_cam
generic map(
G_VSYN_ACTIVE => G_VSYN_ACTIVE
)
port map(
p_in_vd            => p_in_vd,
p_in_vs            => p_in_vin_vs,
p_in_hs            => p_in_vin_hs,
p_in_vclk          => p_in_vin_clk,

p_out_vfr_prm      => i_vfr_prm,

p_out_vbufin_d     => i_vin_dout,--i_vbufin_dout,
p_in_vbufin_rd     => t_vbufin_rd,--i_vbufin_rd,
p_out_vbufin_empty => t_vbufin_empty,--i_vbufin_empty,
p_in_vbufin_rdclk  => g_memclk,

p_in_rst           => i_vctrl_rst
);

t_vbufin_rd<= not t_vbufin_empty;

m_vctrl : cfg2ram_ctrl
generic map(
G_SIM => G_SIM,
G_MEM_AWIDTH => CI_MEM_AWIDTH,
G_MEM_DWIDTH => CI_MEM_DWIDTH
)
port map(
-------------------------------
--
-------------------------------
p_in_rbuf_cfg        => i_hdd_rbuf_cfg,

----------------------------
--����� � ��/��� �������������
----------------------------
--in
p_in_vbufin_d         => i_vbufin_dout,
p_out_vbufin_rd       => i_vbufin_rd,
p_in_vbufin_empty     => i_vbufin_empty,
--out
p_out_vbufout_d       => i_vbufout_din,
p_out_vbufout_wr      => i_vbufout_wr,
p_in_vbufout_full     => i_vbufout_full,

---------------------------------
--����� � mem_ctrl.vhd
---------------------------------
--CH WRITE
p_out_memwr           => i_memch0_in_bank(0), --: out   TMemIN;
p_in_memwr            => i_memch0_out_bank(0),--: in    TMemOUT;
--CH READ
p_out_memrd           => i_memch1_in_bank(0), --: out   TMemIN;
p_in_memrd            => i_memch1_out_bank(0),--: in    TMemOUT;

-------------------------------
--���������������
-------------------------------
p_out_tst             => tst_vctrl_out,

-------------------------------
--System
-------------------------------
p_in_clk              => g_memclk,
p_in_rst              => i_vctrl_rst
);


--***********************************************************
--���������� RAM
--***********************************************************
m_mem_ctrl : mem_ctrl
generic map(
G_SIM => G_SIM
)
port map(
------------------------------------
--User Post
------------------------------------
p_in_memch0     => i_memch0_in_bank, --: in    TMemINBank;
p_out_memch0    => i_memch0_out_bank,--: out   TMemOUTBank;

p_in_memch1     => i_memch1_in_bank, --: in    TMemINBank;
p_out_memch1    => i_memch1_out_bank,--: out   TMemOUTBank;

------------------------------------
--Memory physical interface
------------------------------------
p_out_phymem    => i_phymem_out,
p_inout_phymem  => i_phymem_inout,

------------------------------------
--Memory status
------------------------------------
p_out_mem_rdy   => i_mem_ctrl_rdy,

------------------------------------
--System
------------------------------------
p_out_pll_gclkusr => open,--g_memclk,--300MHz
--c5_rst0         : out   std_logic;
p_in_clk        => g_memclk,--g_hdd_dcm_gclk300M,--
p_in_rst        => i_mem_ctrl_rst
);

p_out_mcb5_a        <= i_phymem_out  (0).a;
p_out_mcb5_ba       <= i_phymem_out  (0).ba;
p_out_mcb5_ras_n    <= i_phymem_out  (0).ras_n;
p_out_mcb5_cas_n    <= i_phymem_out  (0).cas_n;
p_out_mcb5_we_n     <= i_phymem_out  (0).we_n;
p_out_mcb5_odt      <= i_phymem_out  (0).odt;
p_out_mcb5_cke      <= i_phymem_out  (0).cke;
p_out_mcb5_dm       <= i_phymem_out  (0).dm;
p_out_mcb5_udm      <= i_phymem_out  (0).udm;
p_out_mcb5_ck       <= i_phymem_out  (0).ck;
p_out_mcb5_ck_n     <= i_phymem_out  (0).ck_n;
p_inout_mcb5_dq     <= i_phymem_inout(0).dq;
p_inout_mcb5_udqs   <= i_phymem_inout(0).udqs;
p_inout_mcb5_udqs_n <= i_phymem_inout(0).udqs_n;
p_inout_mcb5_dqs    <= i_phymem_inout(0).dqs;
p_inout_mcb5_dqs_n  <= i_phymem_inout(0).dqs_n;
p_inout_mcb5_rzq    <= i_phymem_inout(0).rzq;
p_inout_mcb5_zio    <= i_phymem_inout(0).zio;

p_out_mcb1_a        <= i_phymem_out  (1).a;
p_out_mcb1_ba       <= i_phymem_out  (1).ba;
p_out_mcb1_ras_n    <= i_phymem_out  (1).ras_n;
p_out_mcb1_cas_n    <= i_phymem_out  (1).cas_n;
p_out_mcb1_we_n     <= i_phymem_out  (1).we_n;
p_out_mcb1_odt      <= i_phymem_out  (1).odt;
p_out_mcb1_cke      <= i_phymem_out  (1).cke;
p_out_mcb1_dm       <= i_phymem_out  (1).dm;
p_out_mcb1_udm      <= i_phymem_out  (1).udm;
p_out_mcb1_ck       <= i_phymem_out  (1).ck;
p_out_mcb1_ck_n     <= i_phymem_out  (1).ck_n;
p_inout_mcb1_dq     <= i_phymem_inout(1).dq;
p_inout_mcb1_udqs   <= i_phymem_inout(1).udqs;
p_inout_mcb1_udqs_n <= i_phymem_inout(1).udqs_n;
p_inout_mcb1_dqs    <= i_phymem_inout(1).dqs;
p_inout_mcb1_dqs_n  <= i_phymem_inout(1).dqs_n;
p_inout_mcb1_rzq    <= i_phymem_inout(1).rzq;
p_inout_mcb1_zio    <= i_phymem_inout(1).zio;

--***********************************************************
--������ ���������� - dsn_hdd.vhd
--***********************************************************
gen_sata_gt : for i in 0 to C_SH_COUNT_MAX(C_PCFG_HDD_COUNT-1)-1 generate
  ibufds_hdd_gt_refclk : IBUFDS port map(I  => p_in_sata_clk_p(i), IB => p_in_sata_clk_n(i), O => i_hdd_gt_refclk150(i));
end generate gen_sata_gt;

m_hdd : dsn_hdd
generic map(
G_MODULE_USE=> C_PCFG_HDD_USE,
G_HDD_COUNT => C_PCFG_HDD_COUNT,
G_GT_DBUS   => C_PCFG_HDD_GT_DBUS,
G_DBG       => C_PCFG_HDD_DBG,
G_DBGCS     => C_PCFG_HDD_DBGCS,
G_SIM       => G_SIM
)
port map(
-------------------------------
--���������������� ������ dsn_hdd.vhd (p_in_cfg_clk domain)
-------------------------------
p_in_cfg_if           => C_HDD_CFGIF_UART,
p_in_cfg_clk          => g_sata_refclkout,

p_in_cfg_adr          => i_cfg_adr(7 downto 0),
p_in_cfg_adr_ld       => i_cfg_adr_ld,
p_in_cfg_adr_fifo     => i_cfg_adr_fifo,

p_in_cfg_txdata       => i_cfg_txd,
p_in_cfg_wd           => i_cfg_wd,
p_out_cfg_txrdy       => i_cfg_txrdy,

p_out_cfg_rxdata      => i_cfg_rxd,
p_in_cfg_rd           => i_cfg_rd,
p_out_cfg_rxrdy       => i_cfg_rxrdy,

p_in_cfg_done         => i_cfg_done,
p_in_cfg_rst          => i_sys_rst,

-------------------------------
--STATUS ������ dsn_hdd.vhd
-------------------------------
p_out_hdd_rdy         => i_hdd_module_rdy,
p_out_hdd_error       => i_hdd_module_error,
p_out_hdd_busy        => i_hdd_busy,
p_out_hdd_irq         => open, --i_hdd_hirq,
p_out_hdd_done        => i_hdd_done,

-------------------------------
--����� � �����������/����������� ������ ����������
-------------------------------
p_out_rbuf_cfg        => i_hdd_rbuf_cfg,
p_in_rbuf_status      => i_hdd_rbuf_status,

p_in_hdd_txd          => i_hdd_txdata,
p_in_hdd_txd_wr       => i_hdd_txdata_wd,
p_out_hdd_txbuf_pfull => i_hdd_txbuf_pfull,
p_out_hdd_txbuf_full  => i_hdd_txbuf_full,
p_out_hdd_txbuf_empty => i_hdd_txbuf_empty,

p_out_hdd_rxd         => i_hdd_rxdata,
p_in_hdd_rxd_rd       => i_hdd_rxdata_rd,
p_out_hdd_rxbuf_empty => i_hdd_rxbuf_empty,
p_out_hdd_rxbuf_pempty=> i_hdd_rxbuf_pempty,

-------------------------------
--Sata Driver
-------------------------------
p_out_sata_txn        => p_out_sata_txn,
p_out_sata_txp        => p_out_sata_txp,
p_in_sata_rxn         => p_in_sata_rxn,
p_in_sata_rxp         => p_in_sata_rxp,

p_in_sata_refclk      => i_hdd_gt_refclk150,
p_out_sata_refclkout  => g_sata_refclkout,
p_out_sata_gt_plldet  => i_hdd_gt_plldet,
p_out_sata_dcm_lock   => i_hdd_dcm_lock,
p_out_sata_dcm_gclk2div=> g_hdd_dcm_gclk75M,
p_out_sata_dcm_gclk2x  => g_hdd_dcm_gclk300M,
p_out_sata_dcm_gclk0   => g_hdd_dcm_gclk150M,

-------------------------------
--��������������� ����
-------------------------------
p_in_tst              => (others=>'0'),--i_hdd_tst_in,
p_out_tst             => i_hdd_tst_out,

-------------------------------
--Debug/Sim
-------------------------------
p_out_dbgcs                 => i_hdd_dbgcs,
p_out_dbgled                => i_hdd_dbgled,

p_out_sim_gt_txdata         => open,--i_hdd_sim_gt_txdata,
p_out_sim_gt_txcharisk      => open,--i_hdd_sim_gt_txcharisk,
p_out_sim_gt_txcomstart     => open,--i_hdd_sim_gt_txcomstart,
p_in_sim_gt_rxdata          => i_hdd_sim_gt_rxdata,
p_in_sim_gt_rxcharisk       => i_hdd_sim_gt_rxcharisk,
p_in_sim_gt_rxstatus        => i_hdd_sim_gt_rxstatus,
p_in_sim_gt_rxelecidle      => i_hdd_sim_gt_rxelecidle,
p_in_sim_gt_rxdisperr       => i_hdd_sim_gt_rxdisperr,
p_in_sim_gt_rxnotintable    => i_hdd_sim_gt_rxnotintable,
p_in_sim_gt_rxbyteisaligned => i_hdd_sim_gt_rxbyteisaligned,
p_out_gt_sim_rst            => open,--i_hdd_sim_gt_sim_rst,
p_out_gt_sim_clk            => open,--i_hdd_sim_gt_sim_clk,

-------------------------------
--System
-------------------------------
p_in_clk           => g_sata_refclkout,--p_in_mem_ctrl_clk,--
p_in_rst           => i_hdd_rst
);

gen_satah: for i in 0 to C_HDD_COUNT_MAX-1 generate
i_hdd_sim_gt_rxdata(i)<=(others=>'0');
i_hdd_sim_gt_rxcharisk(i)<=(others=>'0');
i_hdd_sim_gt_rxstatus(i)<=(others=>'0');
i_hdd_sim_gt_rxelecidle(i)<='0';
i_hdd_sim_gt_rxdisperr(i)<=(others=>'0');
i_hdd_sim_gt_rxnotintable(i)<=(others=>'0');
i_hdd_sim_gt_rxbyteisaligned(i)<='0';
end generate gen_satah;

i_hdd_rbuf_status.err<='0';
i_hdd_rbuf_status.err_type.vinbuf_full<='0';
i_hdd_rbuf_status.err_type.rambuf_full<='0';
i_hdd_rbuf_status.done <='0';
i_hdd_rbuf_status.hwlog_size<=(others=>'0');


--***********************************************************
--����� � RAM
--***********************************************************
--RAM<-CFG
m_txram : hdd_ram_hfifo
port map(
din         => i_hdd_rbuf_cfg.ram_wr_i.din,
wr_en       => i_hdd_rbuf_cfg.ram_wr_i.wr,
wr_clk      => i_hdd_rbuf_cfg.ram_wr_i.clk,

dout        => i_hdd_txdata,
rd_en       => i_ram_txbuf_rd,
rd_clk      => g_memclk,--g_sata_refclkout,

full        => i_ram_txbuf_full,
almost_full => i_ram_txbuf_afull,
empty       => i_ram_txbuf_empty,

--clk         => p_in_clk,
rst         => i_ram_reset_buf
);

i_hdd_rbuf_status.ram_wr_o.wr_rdy<= not i_ram_txbuf_afull;
i_hdd_txdata_wd<=(not i_ram_txbuf_empty and not i_hdd_txbuf_pfull) when i_hdd_tst_out(7)='1' else '0';
i_ram_txbuf_rd<=i_hdd_txdata_wd when i_hdd_tst_out(7)='1' else i_vbufin_rd;

i_vbufin_dout<=i_hdd_txdata;
i_vbufin_empty<='1' when i_hdd_tst_out(7)='1' else i_ram_txbuf_empty;


--RAM->CFG
m_rxram : hdd_ram_hfifo
port map(
din         => i_ram_rxbuf_din, --i_hdd_rxdata,
wr_en       => i_ram_rxbuf_wr, --i_hdd_rxdata_rd,
wr_clk      => g_memclk,--g_sata_refclkout,

dout        => i_hdd_rbuf_status.ram_wr_o.dout,
rd_en       => i_hdd_rbuf_cfg.ram_wr_i.rd,
rd_clk      => i_hdd_rbuf_cfg.ram_wr_i.clk,

full        => i_ram_rxbuf_full,
almost_full => i_ram_rxbuf_afull,
empty       => i_ram_rxbuf_empty,

--clk         => p_in_clk,
rst         => i_ram_reset_buf
);

i_hdd_rbuf_status.ram_wr_o.rd_rdy<= not i_ram_rxbuf_afull;
i_hdd_rxdata_rd<=(not i_hdd_rxbuf_empty and not i_ram_rxbuf_afull) when i_hdd_tst_out(7)='1' else '0';
i_ram_rxbuf_wr<=i_hdd_rxdata_rd when i_hdd_tst_out(7)='1' else i_vbufout_wr;
i_ram_rxbuf_din<=i_hdd_rxdata when i_hdd_tst_out(7)='1' else i_vbufout_din;

i_vbufout_full<=i_ram_rxbuf_afull;


--***********************************************************
--��������������� �������
--***********************************************************
m_test01: fpga_test_01
generic map(
G_BLINK_T05   =>10#250#, -- 1/2 ������� ������� ����������.(����� � ms)
G_CLK_T05us   =>10#75#   -- 05us - 150MHz
)
port map(
p_out_test_led => i_test01_led,
p_out_test_done=> open,

p_out_1us      => open,
p_out_1ms      => open,
-------------------------------
--System
-------------------------------
p_in_clk       => g_sata_refclkout,
p_in_rst       => i_sys_rst
);


m_cfgdev : cfgdev_ftdi
port map(
-------------------------------
--����� � FTDI
-------------------------------
p_inout_ftdi_d       => p_inout_ftdi_d,
p_out_ftdi_rd_n      => p_out_ftdi_rd_n,
p_out_ftdi_wr_n      => p_out_ftdi_wr_n,
p_in_ftdi_txe_n      => p_in_ftdi_txe_n,
p_in_ftdi_rxf_n      => p_in_ftdi_rxf_n,
p_in_ftdi_pwren_n    => p_in_ftdi_pwren_n,

-------------------------------
--
-------------------------------
p_out_module_rdy     => open,
p_out_module_error   => open,

-------------------------------
--������/������ ���������������� ���������� ���-��
-------------------------------
p_out_cfg_dadr       => i_dev_adr,
p_out_cfg_radr       => i_cfg_adr,
p_out_cfg_radr_ld    => i_cfg_adr_ld,
p_out_cfg_radr_fifo  => i_cfg_adr_fifo,
p_out_cfg_wr         => i_cfg_wd,
p_out_cfg_rd         => i_cfg_rd,
p_out_cfg_txdata     => i_cfg_txd,
p_in_cfg_rxdata      => i_cfg_rxd,
p_in_cfg_txrdy       => i_cfg_txrdy,
p_in_cfg_rxrdy       => i_cfg_rxrdy,

p_out_cfg_done       => i_cfg_done,
p_in_cfg_clk         => g_sata_refclkout,

-------------------------------
--���������������
-------------------------------
p_in_tst             => (others=>'0'),
p_out_tst            => open,--i_cfg_tstout,

-------------------------------
--System
-------------------------------
p_in_rst => i_sys_rst
);

--i_hdd_tst_in(31 downto 0)<=(others=>'0');

--HDD LEDs:
--SATA0 (�� ����� SATA1)
p_out_led(2)<=i_hdd_dbgled(0).link;
p_out_led(4)<=i_hdd_dbgled(0).rdy;
p_out_TP(0) <=i_hdd_dbgled(0).err and i_test01_led;
p_out_TP(1) <=i_hdd_dbgled(0).busy;

--SATA1 (�� ����� SATA0)
p_out_led(3)<=i_hdd_dbgled(1).link;
p_out_led(5)<=i_hdd_dbgled(1).rdy;
p_out_TP(2) <=i_hdd_dbgled(1).err and i_test01_led;
p_out_TP(3) <=i_hdd_dbgled(1).busy;

--SATA2 (�� ����� SATA3)
p_out_led(0)<=i_mem_ctrl_rdy(0);--i_hdd_dbgled(2).link;
p_out_led(7)<=i_ram_rxbuf_empty;--i_hdd_dbgled(2).rdy;
p_out_TP(6) <=i_hdd_dbgled(2).err and i_test01_led;
p_out_TP(7) <=i_hdd_dbgled(2).busy;

--SATA3 (�� ����� SATA2)
p_out_led(1)<=i_hdd_dbgled(3).link;
p_out_led(6)<=i_hdd_dbgled(3).rdy;
p_out_TP(4) <=i_hdd_dbgled(3).err and i_test01_led;
p_out_TP(5) <=i_hdd_dbgled(3).busy;




--gen_dbgcs : if strcmp(C_PCFG_HDD_DBGCS,"ON") generate
--
----m_dbgcs_icon : dbgcs_iconx3
----port map(
----CONTROL0 => i_dbgcs_sh0_spd,
----CONTROL1 => i_dbgcs_hdd0_layer,
----CONTROL2 => i_dbgcs_hdd1_layer
----);
----
----
------//### HDD0_SPD: ########
----m_dbgcs_sh0_spd : dbgcs_sata_layer
----port map
----(
----CONTROL => i_dbgcs_sh0_spd,
----CLK     => i_hdd_dbgcs.sh(0).spd.clk,
----DATA    => i_hdd_dbgcs.sh(0).spd.data(122 downto 0),
----TRIG0   => i_hdd_dbgcs.sh(0).spd.trig0(41 downto 0)
----);
----
------//### HDD0: ########
----m_dbgcs_hdd0_layer : dbgcs_sata_raid --dbgcs_sata_layer
----port map
----(
----CONTROL => i_dbgcs_hdd0_layer,
----CLK     => i_hdd_dbgcs.sh(0).layer.clk,
----DATA    => i_hdd_dbgcs.sh(0).layer.data(172 downto 0),--(122 downto 0),
----TRIG0   => i_hdd0layer_dbgcs.trig0(41 downto 0)
----);
----
----i_hdd0layer_dbgcs.trig0(19 downto 0)<=i_hdd_dbgcs.sh(0).layer.trig0(19 downto 0);--llayer
----i_hdd0layer_dbgcs.trig0(20)<=i_hdd_dbgcs.sh(0).layer.data(160);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+1);--//C_PSTAT_DET_ESTABLISH_ON_BIT
----i_hdd0layer_dbgcs.trig0(21)<=i_hdd_dbgcs.sh(0).layer.data(161);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+0);--//C_PSTAT_DET_DEV_ON_BIT
----i_hdd0layer_dbgcs.trig0(22)<=i_hdd_dbgcs.sh(0).layer.data(162);--<=p_in_txelecidle;
----i_hdd0layer_dbgcs.trig0(23)<=i_hdd_dbgcs.sh(0).layer.data(163);--<=p_in_rxelecidle;
----i_hdd0layer_dbgcs.trig0(24)<=i_hdd_dbgcs.sh(0).layer.data(164);--<=p_in_txcomstart;
----i_hdd0layer_dbgcs.trig0(25)<=i_hdd_dbgcs.sh(0).layer.data(167);--<=p_in_rxcdrreset;
----i_hdd0layer_dbgcs.trig0(41 downto 26)<=i_hdd_dbgcs.sh(0).layer.trig0(41 downto 26);--llayer
----
------//### HDD1: ########
----gen_hdd1 : if C_PCFG_HDD_COUNT=1 generate
----m_dbgcs_hdd1_layer : dbgcs_sata_raid --dbgcs_sata_layer
----port map
----(
----CONTROL => i_dbgcs_hdd1_layer,
----CLK     => i_hdd_dbgcs.sh(0).layer.clk,
----DATA    => i_hdd_dbgcs.sh(0).layer.data(172 downto 0),--(122 downto 0),
----TRIG0   => i_hdd1layer_dbgcs.trig0(41 downto 0)
----);
----
----i_hdd1layer_dbgcs.trig0(19 downto 0)<=i_hdd_dbgcs.sh(0).layer.trig0(19 downto 0);--llayer
----i_hdd1layer_dbgcs.trig0(20)<=i_hdd_dbgcs.sh(0).layer.data(160);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+1);--//C_PSTAT_DET_ESTABLISH_ON_BIT
----i_hdd1layer_dbgcs.trig0(21)<=i_hdd_dbgcs.sh(0).layer.data(161);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+0);--//C_PSTAT_DET_DEV_ON_BIT
----i_hdd1layer_dbgcs.trig0(22)<=i_hdd_dbgcs.sh(0).layer.data(162);--<=p_in_txelecidle;
----i_hdd1layer_dbgcs.trig0(23)<=i_hdd_dbgcs.sh(0).layer.data(163);--<=p_in_rxelecidle;
----i_hdd1layer_dbgcs.trig0(24)<=i_hdd_dbgcs.sh(0).layer.data(164);--<=p_in_txcomstart;
----i_hdd1layer_dbgcs.trig0(25)<=i_hdd_dbgcs.sh(0).layer.data(167);--<=p_in_rxcdrreset;
----i_hdd1layer_dbgcs.trig0(41 downto 26)<=i_hdd_dbgcs.sh(0).layer.trig0(41 downto 26);--llayer
----end generate gen_hdd1;
----
----gen_hdd2 : if C_PCFG_HDD_COUNT=2 generate
----m_dbgcs_hdd1_layer : dbgcs_sata_raid --dbgcs_sata_layer
----port map
----(
----CONTROL => i_dbgcs_hdd1_layer,
----CLK     => i_hdd_dbgcs.sh(1).layer.clk,
----DATA    => i_hdd_dbgcs.sh(1).layer.data(172 downto 0),--(122 downto 0),
----TRIG0   => i_hdd1layer_dbgcs.trig0(41 downto 0)
----);
----
----i_hdd1layer_dbgcs.trig0(19 downto 0)<=i_hdd_dbgcs.sh(1).layer.trig0(19 downto 0);--llayer
----i_hdd1layer_dbgcs.trig0(20)<=i_hdd_dbgcs.sh(1).layer.data(160);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+1);--//C_PSTAT_DET_ESTABLISH_ON_BIT
----i_hdd1layer_dbgcs.trig0(21)<=i_hdd_dbgcs.sh(1).layer.data(161);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+0);--//C_PSTAT_DET_DEV_ON_BIT
----i_hdd1layer_dbgcs.trig0(22)<=i_hdd_dbgcs.sh(1).layer.data(162);--<=p_in_txelecidle;
----i_hdd1layer_dbgcs.trig0(23)<=i_hdd_dbgcs.sh(1).layer.data(163);--<=p_in_rxelecidle;
----i_hdd1layer_dbgcs.trig0(24)<=i_hdd_dbgcs.sh(1).layer.data(164);--<=p_in_txcomstart;
----i_hdd1layer_dbgcs.trig0(25)<=i_hdd_dbgcs.sh(1).layer.data(167);--<=p_in_rxcdrreset;
----i_hdd1layer_dbgcs.trig0(41 downto 26)<=i_hdd_dbgcs.sh(1).layer.trig0(41 downto 26);--llayer
----end generate gen_hdd2;
----
----gen_hdd3 : if C_PCFG_HDD_COUNT>2 generate
----m_dbgcs_hdd1_layer : dbgcs_sata_raid --dbgcs_sata_layer
----port map
----(
----CONTROL => i_dbgcs_hdd1_layer,
----CLK     => i_hdd_dbgcs.sh(2).layer.clk,
----DATA    => i_hdd_dbgcs.sh(2).layer.data(172 downto 0),--(122 downto 0),
----TRIG0   => i_hdd1layer_dbgcs.trig0(41 downto 0)
----);
----
----i_hdd1layer_dbgcs.trig0(19 downto 0)<=i_hdd_dbgcs.sh(2).layer.trig0(19 downto 0);--llayer
----i_hdd1layer_dbgcs.trig0(20)<=i_hdd_dbgcs.sh(2).layer.data(160);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+1);--//C_PSTAT_DET_ESTABLISH_ON_BIT
----i_hdd1layer_dbgcs.trig0(21)<=i_hdd_dbgcs.sh(2).layer.data(161);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+0);--//C_PSTAT_DET_DEV_ON_BIT
----i_hdd1layer_dbgcs.trig0(22)<=i_hdd_dbgcs.sh(2).layer.data(162);--<=p_in_txelecidle;
----i_hdd1layer_dbgcs.trig0(23)<=i_hdd_dbgcs.sh(2).layer.data(163);--<=p_in_rxelecidle;
----i_hdd1layer_dbgcs.trig0(24)<=i_hdd_dbgcs.sh(2).layer.data(164);--<=p_in_txcomstart;
----i_hdd1layer_dbgcs.trig0(25)<=i_hdd_dbgcs.sh(2).layer.data(167);--<=p_in_rxcdrreset;
----i_hdd1layer_dbgcs.trig0(41 downto 26)<=i_hdd_dbgcs.sh(2).layer.trig0(41 downto 26);--llayer
------
------m_dbgcs_hdd1_layer : dbgcs_sata_raid --dbgcs_sata_layer
------port map
------(
------CONTROL => i_dbgcs_hdd1_layer,
------CLK     => i_hdd_dbgcs.sh(3).layer.clk,
------DATA    => i_hdd_dbgcs.sh(3).layer.data(172 downto 0),--(122 downto 0),
------TRIG0   => i_hdd1layer_dbgcs.trig0(41 downto 0)
------);
------
------i_hdd1layer_dbgcs.trig0(19 downto 0)<=i_hdd_dbgcs.sh(3).layer.trig0(19 downto 0);--llayer
------i_hdd1layer_dbgcs.trig0(20)<=i_hdd_dbgcs.sh(3).layer.data(160);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+1);--//C_PSTAT_DET_ESTABLISH_ON_BIT
------i_hdd1layer_dbgcs.trig0(21)<=i_hdd_dbgcs.sh(3).layer.data(161);--<=p_in_alstatus.sstatus(C_ASSTAT_DET_BIT_L+0);--//C_PSTAT_DET_DEV_ON_BIT
------i_hdd1layer_dbgcs.trig0(22)<=i_hdd_dbgcs.sh(3).layer.data(162);--<=p_in_txelecidle;
------i_hdd1layer_dbgcs.trig0(23)<=i_hdd_dbgcs.sh(3).layer.data(163);--<=p_in_rxelecidle;
------i_hdd1layer_dbgcs.trig0(24)<=i_hdd_dbgcs.sh(3).layer.data(164);--<=p_in_txcomstart;
------i_hdd1layer_dbgcs.trig0(25)<=i_hdd_dbgcs.sh(3).layer.data(167);--<=p_in_rxcdrreset;
------i_hdd1layer_dbgcs.trig0(41 downto 26)<=i_hdd_dbgcs.sh(3).layer.trig0(41 downto 26);--llayer
----end generate gen_hdd3;
--
--
----//### HDD_RAID: ########
--m_dbgcs_icon : dbgcs_iconx1
--port map(
--CONTROL0 => i_dbgcs_hdd_raid
--);
--
--m_dbgcs_sh0_raid : dbgcs_sata_raid
--port map(
--CONTROL => i_dbgcs_hdd_raid,
--CLK     => i_hdd_dbgcs.raid.clk,
--DATA    => i_hddraid_dbgcs.data(172 downto 0),--(122 downto 0),
--TRIG0   => i_hddraid_dbgcs.trig0(41 downto 0)
--);
--
----//-------- TRIG: ------------------
--i_hddraid_dbgcs.trig0(18 downto 0)<=i_hdd_dbgcs.raid.trig0(18 downto 0);
--i_hddraid_dbgcs.trig0(19)<=i_hdd_rbuf_cfg.ram_wr_i.rd;
--
----//SH0
--i_hddraid_dbgcs.trig0(24 downto 20)<=i_hdd_dbgcs.sh(0).layer.trig0(34 downto 30);--llayer
--i_hddraid_dbgcs.trig0(29 downto 25)<=i_hdd_dbgcs.sh(0).layer.trig0(39 downto 35);--tlayer
----//SH1
--i_hddraid_dbgcs.trig0(34 downto 30)<=i_hdd_dbgcs.sh(2).layer.trig0(34 downto 30);--llayer
--i_hddraid_dbgcs.trig0(39 downto 35)<=i_hdd_dbgcs.sh(2).layer.trig0(39 downto 35);--tlayer
--
--i_hddraid_dbgcs.trig0(40)<=i_hdd_txbuf_empty;
--i_hddraid_dbgcs.trig0(41)<=i_hdd_txbuf_pfull;
--
--
----//-------- VIEW: ------------------
--i_hddraid_dbgcs.data(28 downto 0)<=i_hdd_dbgcs.raid.data(28 downto 0);
--i_hddraid_dbgcs.data(29)<=i_hdd_txbuf_pfull;
--
----//SH0
--i_hddraid_dbgcs.data(34 downto 30)<=i_hdd_dbgcs.sh(0).layer.trig0(34 downto 30);--llayer
--i_hddraid_dbgcs.data(39 downto 35)<=i_hdd_dbgcs.sh(0).layer.trig0(39 downto 35);--tlayer
--i_hddraid_dbgcs.data(55 downto 40)<=i_hdd_dbgcs.sh(0).layer.data(65 downto 50);--p_in_ll_rxd(15 downto 0) ---(115 downto 100);--tst_cnt
------i_hddraid_dbgcs.data(55 downto 40)<=i_hdd_dbgcs.sh(0).layer.data(65 downto 50);--p_in_ll_rxd(15 downto 0);--llayer->tlayer
----i_hddraid_dbgcs.data(55 downto 40)<=i_hdd_dbgcs.sh(0).layer.data(97 downto 82);--p_in_ll_txd(15 downto 0);--llayer<-tlayer
--i_hddraid_dbgcs.data(56)          <=i_hdd_dbgcs.sh(0).layer.data(49);--p_in_ll_rxd_wr; --llayer->tlayer
--i_hddraid_dbgcs.data(57)          <=i_hdd_dbgcs.sh(0).layer.data(116);--p_in_ll_txd_rd; --llayer<-tlayer
--i_hddraid_dbgcs.data(58)          <=i_hdd_dbgcs.sh(0).layer.data(118);--<=p_in_dbg.llayer.txbuf_status.aempty; --p_in_gt_txcharisk(0);
--i_hddraid_dbgcs.data(59)          <=i_hdd_dbgcs.sh(0).layer.data(119);--<=p_in_dbg.llayer.txbuf_status.empty; --p_in_gt_txcharisk(1);
--i_hddraid_dbgcs.data(60)          <=i_hdd_dbgcs.sh(0).layer.data(98);--<=p_in_dbg.llayer.rxbuf_status.pfull; --p_in_gt_rxcharisk(0);
--i_hddraid_dbgcs.data(61)          <=i_hdd_dbgcs.sh(0).layer.data(99);--<=p_in_dbg.llayer.txbuf_status.pfull; --p_in_gt_rxcharisk(1);
--i_hddraid_dbgcs.data(62)          <=i_hdd_dbgcs.sh(0).layer.data(117);--<=p_in_dbg.llayer.txd_close;
--
----//SH1
--i_hddraid_dbgcs.data(67 downto 63)<=i_hdd_dbgcs.sh(2).layer.trig0(34 downto 30);--llayer
--i_hddraid_dbgcs.data(72 downto 68)<=i_hdd_dbgcs.sh(2).layer.trig0(39 downto 35);--tlayer
--i_hddraid_dbgcs.data(88 downto 73)<=i_hdd_dbgcs.sh(2).layer.data(65 downto 50);--p_in_ll_rxd(15 downto 0) ---(115 downto 100);--tst_cnt
------i_hddraid_dbgcs.data(88 downto 73)<=i_hdd_dbgcs.sh(2).layer.data(65 downto 50);--p_in_ll_rxd(15 downto 0);--llayer->tlayer
----i_hddraid_dbgcs.data(88 downto 73)<=i_hdd_dbgcs.sh(2).layer.data(97 downto 82);--p_in_ll_txd(15 downto 0);--llayer<-tlayer
--i_hddraid_dbgcs.data(89)          <=i_hdd_dbgcs.sh(2).layer.data(49);--p_in_ll_rxd_wr; --llayer->tlayer
--i_hddraid_dbgcs.data(90)          <=i_hdd_dbgcs.sh(2).layer.data(116);--p_in_ll_txd_rd; --llayer<-tlayer
--i_hddraid_dbgcs.data(91)          <=i_hdd_dbgcs.sh(2).layer.data(118);--<=p_in_dbg.llayer.txbuf_status.aempty; --p_in_gt_txcharisk(0);
--i_hddraid_dbgcs.data(92)          <=i_hdd_dbgcs.sh(2).layer.data(119);--<=p_in_dbg.llayer.txbuf_status.empty; --p_in_gt_txcharisk(1);
--i_hddraid_dbgcs.data(93)          <=i_hdd_dbgcs.sh(2).layer.data(98);--<=p_in_dbg.llayer.rxbuf_status.pfull; --p_in_gt_rxcharisk(0);
--i_hddraid_dbgcs.data(94)          <=i_hdd_dbgcs.sh(2).layer.data(99);--<=p_in_dbg.llayer.txbuf_status.pfull; --p_in_gt_rxcharisk(1);
--i_hddraid_dbgcs.data(95)          <=i_hdd_done;--i_hdd_rambuf_dbgcs.data(3);--i_hdd_dbgcs.sh(1).layer.data(117);--<=p_in_dbg.llayer.txd_close;
--
----//RAMBUF
--i_hddraid_dbgcs.data(103 downto 100)<=(others=>'0');
--i_hddraid_dbgcs.data(104)<=i_hdd_txbuf_empty;
--i_hddraid_dbgcs.data(105)<=i_hdd_rxbuf_empty;
--i_hddraid_dbgcs.data(106)<=i_hdd_txdata_wd;--RAM->HDD
--i_hddraid_dbgcs.data(107)<=i_hdd_rxdata_rd;--RAM<-HDD
--i_hddraid_dbgcs.data(108)<=i_ram_rxbuf_empty;
--i_hddraid_dbgcs.data(140 downto 109)<=i_hdd_dbgcs.raid.data(161 downto 130);--i_usr_rxd;--RAM<-HDD
--i_hddraid_dbgcs.data(172 downto 141)<=i_hdd_rxdata(31 downto 0);--RAM<-HDD
--
--
--end generate gen_dbgcs;
--
--

--m_dbgcs_icon : dbgcs_iconx2
--port map(
--CONTROL0 => i_dbgcs_hdd_raid,
--CONTROL1 => i_dbgcs_cfg
--);
m_dbgcs_icon : dbgcs_iconx1
port map(
CONTROL0 => i_dbgcs_hdd_raid
);

m_dbgcs_sh0_raid : dbgcs_sata_raid
port map(
CONTROL => i_dbgcs_hdd_raid,
CLK     => g_memclk,--i_hdd_dbgcs.raid.clk,
DATA    => i_hddraid_dbgcs.data(172 downto 0),--(122 downto 0),
TRIG0   => i_hddraid_dbgcs.trig0(41 downto 0)
);

--//-------- TRIG: ------------------
i_hddraid_dbgcs.trig0(0)            <=tst_vctrl_out(0);         --vwriter(0)<=p_in_cfg_mem_start;
i_hddraid_dbgcs.trig0(1)            <=tst_vctrl_out(1);         --vwriter(1)<=i_mem_done;
i_hddraid_dbgcs.trig0(4 downto 2)   <=tst_vctrl_out(4 downto 2);--vwriter(4 downto 2)<=tst_fsm_cs;
i_hddraid_dbgcs.trig0(5)            <=tst_vctrl_out(5);         --vreader(0)<=p_in_cfg_mem_start;
i_hddraid_dbgcs.trig0(6)            <=tst_vctrl_out(6);         --vreader(1)<=i_mem_done;
i_hddraid_dbgcs.trig0(9 downto 7)   <=tst_vctrl_out(9 downto 7);--vreader(4 downto 2)<=tst_fsm_cs;
i_hddraid_dbgcs.trig0(10)           <=tst_vctrl_out(14)        ;--  <=i_vwr_fr_rdy(0);
i_hddraid_dbgcs.trig0(11)           <=tst_vctrl_out(15)        ;--  <=i_vrd_hold(0);
i_hddraid_dbgcs.trig0(12)           <=p_in_vin_vs;--   : in   std_logic;
i_hddraid_dbgcs.trig0(13)           <=p_in_vin_hs;--   : in   std_logic;
i_hddraid_dbgcs.trig0(14)           <=p_in_vout_vs;--   : in   std_logic;
i_hddraid_dbgcs.trig0(15)           <=p_in_vout_hs;--   : in   std_logic;

i_hddraid_dbgcs.trig0(16)           <=i_memch0_in_bank(0).cmd_wr;-- : std_logic;
i_hddraid_dbgcs.trig0(17)           <=i_memch1_in_bank(0).cmd_wr;-- : std_logic;
i_hddraid_dbgcs.trig0(18)           <=tst_syn;
i_hddraid_dbgcs.trig0(19)           <=i_ram_txbuf_rd;--i_ram_txbuf_empty;
i_hddraid_dbgcs.trig0(20)           <=i_ram_rxbuf_wr;--i_ram_rxbuf_empty;


--//-------- VIEW: ------------------
i_hddraid_dbgcs.data(0)             <=tst_vctrl_out(0);         --vwriter(0)<=p_in_cfg_mem_start;
i_hddraid_dbgcs.data(1)             <=tst_vctrl_out(1);         --vwriter(1)<=i_mem_done;
i_hddraid_dbgcs.data(4 downto 2)    <=tst_vctrl_out(4 downto 2);--vwriter(4 downto 2)<=tst_fsm_cs;
i_hddraid_dbgcs.data(5)             <=tst_vctrl_out(5);         --vreader(0)<=p_in_cfg_mem_start;
i_hddraid_dbgcs.data(6)             <=tst_vctrl_out(6);         --vreader(1)<=i_mem_done;
i_hddraid_dbgcs.data(9 downto 7)    <=tst_vctrl_out(9 downto 7);--vreader(4 downto 2)<=tst_fsm_cs;
i_hddraid_dbgcs.data(10)            <=tst_vctrl_out(14)        ;--  <=i_vwr_fr_rdy(0);/ram_start
i_hddraid_dbgcs.data(11)            <=tst_vctrl_out(15)        ;--  <=i_vrd_hold(0);
i_hddraid_dbgcs.data(13 downto 12)  <=tst_vctrl_out(11 downto 10);--<=i_vbuf_wr(0);
i_hddraid_dbgcs.data(15 downto 14)  <=tst_vctrl_out(13 downto 12);--<=i_vbuf_rd(0);
i_hddraid_dbgcs.data(16)            <=i_vbufin_empty;
i_hddraid_dbgcs.data(17)            <=i_vbufout_full;
i_hddraid_dbgcs.data(18)            <=tst_vin_vs; --   : in   std_logic;
i_hddraid_dbgcs.data(19)            <=tst_vin_hs; --   : in   std_logic;
i_hddraid_dbgcs.data(20)            <=tst_vout_vs;--   : in   std_logic;
i_hddraid_dbgcs.data(21)            <=tst_vout_hs;--   : in   std_logic;

i_hddraid_dbgcs.data(27 downto 22)  <=i_memch0_in_bank (0).cmd_bl       ;--: std_logic_vector(5 downto 0);
i_hddraid_dbgcs.data(28)            <=i_memch0_in_bank (0).cmd_wr       ;--: std_logic;
i_hddraid_dbgcs.data(29)            <=i_memch0_out_bank(0).cmdbuf_full  ;--: std_logic;
i_hddraid_dbgcs.data(30)            <=i_memch0_out_bank(0).cmdbuf_empty ;--: std_logic;
i_hddraid_dbgcs.data(31)            <=i_memch0_in_bank (0).txd_wr       ;--: std_logic;
i_hddraid_dbgcs.data(32)            <=i_memch0_out_bank(0).txbuf_full   ;--: std_logic;
i_hddraid_dbgcs.data(33)            <=i_memch0_out_bank(0).txbuf_empty  ;--: std_logic;
i_hddraid_dbgcs.data(40 downto 34)  <=i_memch0_out_bank(0).txbuf_wrcount;--: std_logic_vector(6 downto 0);
i_hddraid_dbgcs.data(46 downto 41)  <=i_memch1_in_bank (0).cmd_bl       ;--: std_logic_vector(5 downto 0);
i_hddraid_dbgcs.data(47)            <=i_memch1_in_bank (0).cmd_wr       ;--: std_logic;
i_hddraid_dbgcs.data(48)            <=i_memch1_out_bank(0).cmdbuf_full  ;--: std_logic;
i_hddraid_dbgcs.data(49)            <=i_memch1_out_bank(0).cmdbuf_empty ;--: std_logic;
i_hddraid_dbgcs.data(50)            <=i_memch1_in_bank (0).rxd_rd       ;--: std_logic;
i_hddraid_dbgcs.data(51)            <=i_memch1_out_bank(0).rxbuf_full   ;--: std_logic;
i_hddraid_dbgcs.data(52)            <=i_memch1_out_bank(0).rxbuf_empty  ;--: std_logic;
i_hddraid_dbgcs.data(59 downto 53)  <=i_memch1_out_bank(0).rxbuf_rdcount;--: std_logic_vector(6 downto 0);

i_hddraid_dbgcs.data(60)            <=i_ram_txbuf_empty;
i_hddraid_dbgcs.data(61)            <=i_ram_rxbuf_empty;
i_hddraid_dbgcs.data(62)            <=i_vctrl_rst;
i_hddraid_dbgcs.data(63)            <=tst_syn;

i_hddraid_dbgcs.data(95 downto 64)  <=i_vin_dout;--(others=>'0');
i_hddraid_dbgcs.data(96)            <=tst_vctrl_out(16);--<=tst_vwr_out(5);--<=i_mem_cmden;
i_hddraid_dbgcs.data(97)            <=tst_vctrl_out(17);--<=tst_vrd_out(5);--<=i_mem_cmden;
i_hddraid_dbgcs.data(98)            <='0';--tst_vctrl_out(18);--<=tst_vwr_out(6);--<=i_mem_trn_work;
i_hddraid_dbgcs.data(99)            <='0';--tst_vctrl_out(19);--<=tst_vrd_out(6);--<=i_mem_trn_work;

i_hddraid_dbgcs.data(131 downto 100) <=i_hdd_txdata;--Tx --i_memch0_in_bank(0).txd(31 downto 0) ;--i_vbufin_dout
i_hddraid_dbgcs.data(163 downto 132) <=i_ram_rxbuf_din;--i_memch1_out_bank(0).rxd(31 downto 0);--i_vbufout_din;--Rx

i_hddraid_dbgcs.data(164)            <=i_ram_rxbuf_wr;
i_hddraid_dbgcs.data(165)            <=i_ram_txbuf_rd;
i_hddraid_dbgcs.data(166)            <=t_vbufin_rd;



process(g_memclk)
begin
  if g_memclk'event and g_memclk='1' then
    sr_vctrl_rst(0)<=i_vctrl_rst;
    sr_vctrl_rst(1)<=sr_vctrl_rst(0);
    tst_syn<=not sr_vctrl_rst(0) and sr_vctrl_rst(1);

    tst_vin_vs <=p_in_vin_vs ;--   : in   std_logic;
    tst_vin_hs <=p_in_vin_hs ;--   : in   std_logic;
    tst_vout_vs<=p_in_vout_vs;--   : in   std_logic;
    tst_vout_hs<=p_in_vout_hs;--   : in   std_logic;
  end if;
end process;



--m_dbgcs_cfg : dbgcs_sata_raid
--port map(
--CONTROL => i_dbgcs_cfg,
--CLK     => i_hdd_rbuf_cfg.ram_wr_i.clk,--i_hdd_dbgcs.raid.clk,
--DATA    => i_cfg_dbgcs.data(172 downto 0),--(122 downto 0),
--TRIG0   => i_cfg_dbgcs.trig0(41 downto 0)
--);
--
----//-------- TRIG: ------------------
--i_cfg_dbgcs.trig0(0)             <=i_cfg_adr_ld   ;
--i_cfg_dbgcs.trig0(1)             <=i_cfg_adr_fifo ;
--i_cfg_dbgcs.trig0(2)             <=i_cfg_wd       ;
--i_cfg_dbgcs.trig0(5)             <=i_cfg_rd       ;
--i_cfg_dbgcs.trig0(6)             <=i_cfg_txrdy    ;
--i_cfg_dbgcs.trig0(7)             <=i_cfg_rxrdy    ;
--i_cfg_dbgcs.trig0(13 downto 8)   <=i_cfg_adr(5 downto 0);
--i_cfg_dbgcs.trig0(14)            <='0';
--i_cfg_dbgcs.trig0(15)            <='0';
--i_cfg_dbgcs.trig0(16)            <=i_ram_txbuf_empty;
--i_cfg_dbgcs.trig0(17)            <=i_ram_rxbuf_empty;
--
--
----//-------- VIEW: ------------------
--i_cfg_dbgcs.data(0)             <=i_cfg_adr_ld   ;
--i_cfg_dbgcs.data(1)             <=i_cfg_adr_fifo ;
--i_cfg_dbgcs.data(2)             <=i_cfg_wd       ;
--i_cfg_dbgcs.data(5)             <=i_cfg_rd       ;
--i_cfg_dbgcs.data(6)             <=i_cfg_txrdy    ;
--i_cfg_dbgcs.data(7)             <=i_cfg_rxrdy    ;
--i_cfg_dbgcs.data(13 downto 8)   <=i_cfg_adr(5 downto 0);
--
--i_cfg_dbgcs.data(14)            <=i_hdd_tst_out(8);--<=i_ram_d_wcnt;
--i_cfg_dbgcs.data(15)            <='0';
--
--i_cfg_dbgcs.data(31 downto 16)  <=i_cfg_txd;
--i_cfg_dbgcs.data(47 downto 32)  <=i_cfg_rxd;
--
--i_cfg_dbgcs.data(48)            <=i_hdd_rbuf_cfg.ram_wr_i.wr;
--i_cfg_dbgcs.data(49)            <=i_ram_txbuf_empty;
--i_cfg_dbgcs.data(50)            <=i_ram_txbuf_afull;
--
--i_cfg_dbgcs.data(51)            <=i_hdd_rbuf_cfg.ram_wr_i.rd;
--i_cfg_dbgcs.data(52)            <=i_ram_rxbuf_empty;
--i_cfg_dbgcs.data(53)            <=i_ram_rxbuf_afull;
--
--i_cfg_dbgcs.data(63 downto 54)  <=(others=>'0');
--
--i_cfg_dbgcs.data(95 downto 64)  <=i_hdd_rbuf_status.ram_wr_o.dout;
--
--i_cfg_dbgcs.data(172 downto 96) <=(others=>'0');





--END MAIN
end architecture;
