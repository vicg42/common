-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 29.03.2012 13:12:10
-- Module Name : mem_ctrl
--
-- ����������/�������� :
--
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.ext;

library unisim;
use unisim.vcomponents.all;

library work;
use work.mem_ctrl_pkg.all;
use work.mem_wr_pkg.all;

entity mem_ctrl is
generic(
G_SIM : string:= "OFF"
);
port(
------------------------------------
--User Post
------------------------------------
p_in_mem       : in    TMemINBank;
p_out_mem      : out   TMemOUTBank;

------------------------------------
--Memory physical interface
------------------------------------
p_out_phymem   : out   TMEMCTRL_phy_outs;
p_inout_phymem : inout TMEMCTRL_phy_inouts;

------------------------------------
--Memory status
------------------------------------
p_out_status   : out   TMEMCTRL_status;

------------------------------------
--System
------------------------------------
p_out_sys      : out   TMEMCTRL_sysout;
p_in_sys       : in    TMEMCTRL_sysin
);
end;

architecture synth of mem_ctrl is

type TSAXI_ID_t is array (0 to C_MEM_BANK_COUNT-1) of std_logic_vector(C_AXIM_IDWIDTH-1 downto 0);
signal i_saxi_bid      : TSAXI_ID_t;
signal i_saxi_rid      : TSAXI_ID_t;
signal i_clk           : std_logic_vector(C_MEM_BANK_COUNT-1 downto 0);


--MAIN
begin

p_out_sys.clk <= i_clk(0);

gen_bank : for i in 0 to C_MEM_BANK_COUNT-1 generate

p_out_mem(i).axiw.rid <= EXT(i_saxi_bid(i), p_out_mem(i).axiw.rid'length);
p_out_mem(i).axir.rid <= EXT(i_saxi_rid(i), p_out_mem(i).axir.rid'length);
p_out_mem(i).clk <= i_clk(i);

m_mem_core : mem_ctrl_core_axi
port map(
s_axi_aresetn => p_out_mem(i).rstn,
s_axi_clk     => i_clk(i),

-- AXI Slave Interface:
-- Write Address Ports
s_axi_awid     => p_in_mem (i).axiw.aid(C_AXIM_IDWIDTH-1 downto 0),
s_axi_awaddr   => p_in_mem (i).axiw.adr(C_AXI_AWIDTH-1 downto 0)  ,
s_axi_awlen    => p_in_mem (i).axiw.trnlen                        ,
s_axi_awsize   => p_in_mem (i).axiw.dbus                          ,
s_axi_awburst  => p_in_mem (i).axiw.burst                         ,
s_axi_awlock   => p_in_mem (i).axiw.lock                          ,
s_axi_awcache  => p_in_mem (i).axiw.cache                         ,
s_axi_awprot   => p_in_mem (i).axiw.prot                          ,
s_axi_awqos    => p_in_mem (i).axiw.qos                           ,
s_axi_awvalid  => p_in_mem (i).axiw.avalid                        ,
s_axi_awready  => p_out_mem(i).axiw.aready                        ,
-- Write Data Ports
s_axi_wdata    => p_in_mem (i).axiw.data(C_AXIM_DWIDTH-1 downto 0) ,
s_axi_wstrb    => p_in_mem (i).axiw.dbe(C_AXIM_DWIDTH/8-1 downto 0),
s_axi_wlast    => p_in_mem (i).axiw.dlast                         ,
s_axi_wvalid   => p_in_mem (i).axiw.dvalid                        ,
s_axi_wready   => p_out_mem(i).axiw.wready                        ,
-- Write Response Ports
s_axi_bid      => i_saxi_bid(i)(C_AXIM_IDWIDTH-1 downto 0)        ,
s_axi_bresp    => p_out_mem(i).axiw.resp                          ,
s_axi_bvalid   => p_out_mem(i).axiw.rvalid                        ,
s_axi_bready   => p_in_mem (i).axiw.rready                        ,
-- Read Address Ports
s_axi_arid     => p_in_mem (i).axir.aid(C_AXIM_IDWIDTH-1 downto 0),
s_axi_araddr   => p_in_mem (i).axir.adr(C_AXI_AWIDTH-1 downto 0)  ,
s_axi_arlen    => p_in_mem (i).axir.trnlen                        ,
s_axi_arsize   => p_in_mem (i).axir.dbus                          ,
s_axi_arburst  => p_in_mem (i).axir.burst                         ,
s_axi_arlock   => p_in_mem (i).axir.lock                          ,
s_axi_arcache  => p_in_mem (i).axir.cache                         ,
s_axi_arprot   => p_in_mem (i).axir.prot                          ,
s_axi_arqos    => p_in_mem (i).axir.qos                           ,
s_axi_arvalid  => p_in_mem (i).axir.avalid                        ,
s_axi_arready  => p_out_mem(i).axir.aready                        ,
-- Read Data Ports
s_axi_rid      => i_saxi_rid(i)(C_AXIM_IDWIDTH-1 downto 0)        ,
s_axi_rdata    => p_out_mem(i).axir.data(C_AXIM_DWIDTH-1 downto 0) ,
s_axi_rresp    => p_out_mem(i).axir.resp                          ,
s_axi_rlast    => p_out_mem(i).axir.dlast                         ,
s_axi_rvalid   => p_out_mem(i).axir.dvalid                        ,
s_axi_rready   => p_in_mem (i).axir.rready                        ,

--AXI CTRL port
s_axi_ctrl_awvalid => '0',
s_axi_ctrl_awready => open,
s_axi_ctrl_awaddr  => (others=>'0'),
s_axi_ctrl_wvalid  => '0',
s_axi_ctrl_wready  => open,
s_axi_ctrl_wdata   => (others=>'0'),
s_axi_ctrl_bvalid  => open,
s_axi_ctrl_bready  => '1',
s_axi_ctrl_bresp   => open,
s_axi_ctrl_arvalid => '0',
s_axi_ctrl_arready => open,
s_axi_ctrl_araddr  => (others=>'0'),
s_axi_ctrl_rvalid  => open,
s_axi_ctrl_rready  => '1',
s_axi_ctrl_rdata   => open,
s_axi_ctrl_rresp   => open,


-- DDR3 Physical Interface
ddr3_dq         => p_inout_phymem(i).dq   ,
ddr3_addr       => p_out_phymem  (i).a    ,
ddr3_ba         => p_out_phymem  (i).ba   ,
ddr3_ras_n      => p_out_phymem  (i).ras_n,
ddr3_cas_n      => p_out_phymem  (i).cas_n,
ddr3_we_n       => p_out_phymem  (i).we_n ,
ddr3_reset_n    => p_out_phymem  (i).rst_n,
ddr3_cs_n       => p_out_phymem  (i).cs_n ,
ddr3_odt        => p_out_phymem  (i).odt  ,
ddr3_cke        => p_out_phymem  (i).cke  ,
ddr3_dm         => p_out_phymem  (i).dm   ,
ddr3_dqs_p      => p_inout_phymem(i).dqs_p,
ddr3_dqs_n      => p_inout_phymem(i).dqs_n,
ddr3_ck_p       => p_out_phymem  (i).ck_p ,
ddr3_ck_n       => p_out_phymem  (i).ck_n ,

interrupt       => open,

mmcm_locked     => open,

app_sr_req      => '0',
app_sr_active   => open,
app_ref_req     => '0',
app_ref_ack     => open,
app_zq_req      => '0',
app_zq_ack      => open,

device_temp_i   => (others=>'0'),

app_ecc_multiple_err => open,

--Status
init_calib_complete => p_out_status.rdy(i),

--System
sys_clk_i       => p_in_sys.clk    ,
clk_ref_i       => p_in_sys.ref_clk,
sys_rst         => p_in_sys.rst
);

end generate gen_bank;


--END MAIN
end;

