-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 10/26/2007
-- Module Name : prj_def
--
-- Description :
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------
library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;

library work;
use work.vicg_common_pkg.all;
use work.prj_cfg.all;

package prj_def is

--������ �������� FPGA
constant C_FPGA_FIRMWARE_VERSION : integer:=16#0401#;

--//VCTRL
constant C_VIDEO_PKT_HEADER_SIZE : integer:=5;--DWORD

--//HOST
constant C_HDEV_DWIDTH           : integer:=32;--���� ������ p_out_dev_din/p_in_dev_dout ������ dsn_host.vhd

--//--------------------------------------------------------------
--//�������� ������ dsn_host.vhd: (max count HREG - 0x1F)
--//--------------------------------------------------------------
constant C_HREG_FIRMWARE                      : integer:=16#00#;--������ �������� FPGA
constant C_HREG_CTRL                          : integer:=16#01#;--���������� ����������
constant C_HREG_DMAPRM_ADR                    : integer:=16#02#;--����� ������ ���������� � ������ PC ��������� PCI-Express
constant C_HREG_DMAPRM_LEN                    : integer:=16#03#;--������ ������(� ������) ���������� � ������ PC ��������� PCI-Express
constant C_HREG_DEV_CTRL                      : integer:=16#04#;--���������� ����-���� ������������� � ������ dsn_host.vhd
constant C_HREG_DEV_STATUS                    : integer:=16#05#;--������� ��������� ������������ � ������ dsn_host.vhd
constant C_HREG_DEV_DATA                      : integer:=16#06#;--������� ������/������ ������ ����� �� PCIE_DMA
constant C_HREG_IRQ                           : integer:=16#07#;--����������: ���������� + �������
constant C_HREG_MEM_ADR                       : integer:=16#08#;--����� ��� ������������� � FPGA
constant C_HREG_MEM_CTRL                      : integer:=16#09#;
constant C_HREG_VCTRL_FRMRK                   : integer:=16#0A#;--������ ���������� ����������
constant C_HREG_VCTRL_FRERR                   : integer:=16#0B#;
constant C_HREG_TIME                          : integer:=16#0C#;--[31]-overday, [30:26]-����, [25:20]-������, [19:14]-�������, [13:4]-��, [3:0]-����� ���.
constant C_HREG_PCIE                          : integer:=16#0D#;--��� + ������("������" ���������) PCI-Express
constant C_HREG_FUNC                          : integer:=16#0E#;--������������ ������ ������� FPGA
constant C_HREG_FUNCPRM                       : integer:=16#0F#;--���������� � �������
--constant C_HREG_RESERV                        : integer:=...
constant C_HREG_TST0                          : integer:=16#1C#;--�������� ��������
constant C_HREG_TST1                          : integer:=16#1D#;
constant C_HREG_TST2                          : integer:=16#1E#;


--//Register C_HREG_FIRMWARE / Bit Map:
constant C_HREG_FRMWARE_LAST_BIT              : integer:=15;


--//Register C_HREG_CTRL / Bit Map:
constant C_HREG_CTRL_RST_ALL_BIT              : integer:=0;
constant C_HREG_CTRL_RST_MEM_BIT              : integer:=1;
constant C_HREG_CTRL_RST_ETH_BIT              : integer:=2;
constant C_HREG_CTRL_RDDONE_VCTRL_BIT         : integer:=3;
constant C_HREG_CTRL_RST_PULT_BIT             : integer:=4;
constant C_HREG_CTRL_RST_EDEV_BIT             : integer:=5;
constant C_HREG_CTRL_ESYNC_IEDGE_BIT          : integer:=6; --����������� ������ ������ ������� ������������� (0-rise)
constant C_HREG_CTRL_ESYNC_OEDGE_BIT          : integer:=7; --����������� ������ ������� �� ������� ������������� (0-rise)
constant C_HREG_CTRL_ESYNC_MODE_L_BIT         : integer:=8; --'10'-�������, '01'-PPS, '11','00'-���������� �������������
constant C_HREG_CTRL_ESYNC_MODE_M_BIT         : integer:=9; --
constant C_HREG_CTRL_TIME_MODE_BIT            : integer:=10;--��������� ����� (0-����� � �������, 1-�� ������� �������)
constant C_HREG_CTRL_TIME_EN_BIT              : integer:=11;--���������� ������ ����� (1-���������)
constant C_HREG_CTRL_RST_BUP_BIT              : integer:=12;
constant C_HREG_CTRL_RST_VIZIR_BIT            : integer:=13;
constant C_HREG_CTRL_BITCLK_VIZIR_BIT         : integer:=14;--1/0  = bitclk 1MHz/ bitclk 250kHz
constant C_HREG_CTRL_RST_PROM_BIT             : integer:=15;
constant C_HREG_CTRL_EN_SYN120_BUP_BIT        : integer:=16;--���������� ������ � BUP �� ������� 120 ��
                                                            --������������ � PPS GPS (������ 120�� ������� �� ������ m_sync)
constant C_HREG_CTRL_LAST_BIT                 : integer:=C_HREG_CTRL_EN_SYN120_BUP_BIT;


--//Register C_HREG_DEV_CTRL / Bit Map:
constant C_HREG_DEV_CTRL_DRDY_BIT             : integer:=0;
constant C_HREG_DEV_CTRL_DMA_START_BIT        : integer:=1; --(�������� �����)������ ������� ��������
constant C_HREG_DEV_CTRL_DMA_DIR_BIT          : integer:=2; --1/0 � ������/������ ������ ����������������� ����������
constant C_HREG_DEV_CTRL_DMABUF_L_BIT         : integer:=3; --��������� ����� ������ � ����������� PCIE_DMA
constant C_HREG_DEV_CTRL_DMABUF_M_BIT         : integer:=10;
constant C_HREG_DEV_CTRL_DMABUF_COUNT_L_BIT   : integer:=11;--����� ���-�� ������� � ����������� PCIE_DMA
constant C_HREG_DEV_CTRL_DMABUF_COUNT_M_BIT   : integer:=18;
constant C_HREG_DEV_CTRL_ADR_L_BIT            : integer:=19;--����� ����������������� ����������:(C_HDEV_xxx)
constant C_HREG_DEV_CTRL_ADR_M_BIT            : integer:=22;
constant C_HREG_DEV_CTRL_VCH_L_BIT            : integer:=23;--����� ����� ������
constant C_HREG_DEV_CTRL_VCH_M_BIT            : integer:=25;
constant C_HREG_DEV_CTRL_LAST_BIT             : integer:=C_HREG_DEV_CTRL_VCH_M_BIT;--Max 31

--//���� C_HREG_DEV_CTRL_ADR - ������ ���������������� ���������:
constant C_HDEV_CFG_DBUF                      : integer:=0;--������ RX/TX CFG
constant C_HDEV_ETH_DBUF                      : integer:=1;--������ RX/TX ETH
constant C_HDEV_MEM_DBUF                      : integer:=2;--���
constant C_HDEV_VCH_DBUF                      : integer:=3;--����� ���������������
constant C_HDEV_EDEV_DBUF                     : integer:=4;--External Device (������, ���������...)
constant C_HDEV_PULT_DBUF                     : integer:=5;--
constant C_HDEV_VIZIR_DBUF                    : integer:=6;--
constant C_HDEV_BUP_DBUF                      : integer:=7;--���� ���������� ���������
constant C_HDEV_PROM                          : integer:=8;--Bootloader FPGA firmware
constant C_HDEV_COUNT                         : integer:=C_HDEV_PROM+1;
constant C_HDEV_COUNT_MAX                     : integer:=pwr(2, (C_HREG_DEV_CTRL_ADR_M_BIT-C_HREG_DEV_CTRL_ADR_L_BIT+1));

--//Register C_HOST_REG_STATUS_DEV / Bit Map:
--constant RESERV                             : integer:=0;
constant C_HREG_DEV_STATUS_PROM_TXRDY_BIT     : integer:=1;
constant C_HREG_DEV_STATUS_PROM_RXRDY_BIT     : integer:=2;
constant C_HREG_DEV_STATUS_PROM_ERR_BIT       : integer:=3;
constant C_HREG_DEV_STATUS_DMA_BUSY_BIT       : integer:=4; --PCIE_DMA
constant C_HREG_DEV_STATUS_CFG_RDY_BIT        : integer:=5;
constant C_HREG_DEV_STATUS_CFG_RXRDY_BIT      : integer:=6;
constant C_HREG_DEV_STATUS_CFG_TXRDY_BIT      : integer:=7;
constant C_HREG_DEV_STATUS_ETH_RDY_BIT        : integer:=8;
constant C_HREG_DEV_STATUS_ETH_LINK_BIT       : integer:=9;
constant C_HREG_DEV_STATUS_ETH_RXRDY_BIT      : integer:=10;
constant C_HREG_DEV_STATUS_ETH_TXRDY_BIT      : integer:=11;
constant C_HREG_DEV_STATUS_MEMCTRL_RDY_BIT    : integer:=12;
constant C_HREG_DEV_STATUS_EDEV_TXRDY_BIT     : integer:=13;
constant C_HREG_DEV_STATUS_EDEV_RXRDY_BIT     : integer:=14;
constant C_HREG_DEV_STATUS_EDEV_RXERR_BIT     : integer:=15;
constant C_HREG_DEV_STATUS_VCH0_FRRDY_BIT     : integer:=16;
constant C_HREG_DEV_STATUS_VCH1_FRRDY_BIT     : integer:=17;
constant C_HREG_DEV_STATUS_VCH2_FRRDY_BIT     : integer:=18;
constant C_HREG_DEV_STATUS_VCH3_FRRDY_BIT     : integer:=19;
constant C_HREG_DEV_STATUS_VCH4_FRRDY_BIT     : integer:=20;
constant C_HREG_DEV_STATUS_VCH5_FRRDY_BIT     : integer:=21;
constant C_HREG_DEV_STATUS_PULT_TXRDY_BIT     : integer:=22;
constant C_HREG_DEV_STATUS_PULT_RXRDY_BIT     : integer:=23;
constant C_HREG_DEV_STATUS_VIZIR_TXRDY_BIT    : integer:=24;
constant C_HREG_DEV_STATUS_VIZIR_RXRDY_BIT    : integer:=25;
constant C_HREG_DEV_STATUS_VIZIR_RXERR_BIT    : integer:=26;
constant C_HREG_DEV_STATUS_BUP_TXRDY_BIT      : integer:=27;
constant C_HREG_DEV_STATUS_BUP_RXRDY_BIT      : integer:=28;
constant C_HREG_DEV_STATUS_BUP_RXERR_BIT      : integer:=29;
constant C_HREG_DEV_STATUS_LAST_BIT           : integer:=C_HREG_DEV_STATUS_BUP_RXERR_BIT;


--//Register C_HREG_IRQ / Bit Map:
constant C_HREG_IRQ_NUM_L_WBIT                : integer:=0; --����� ��������� ����������
constant C_HREG_IRQ_NUM_M_WBIT                : integer:=4; --
constant C_HREG_IRQ_EN_WBIT                   : integer:=13;--���������� ���������� �� ���������������� ���������
constant C_HREG_IRQ_DIS_WBIT                  : integer:=14;--��������� ���������� �� ���������������� ���������
constant C_HREG_IRQ_CLR_WBIT                  : integer:=15;--����� ������� ���������� �����. ��������� ����������
constant C_HREG_IRQ_LAST_WBIT                 : integer:=C_HREG_IRQ_CLR_WBIT;

constant C_HREG_IRQ_STATUS_L_RBIT             : integer:=0; --������� ���������� ���������� �� �����. ���������
constant C_HREG_IRQ_STATUS_M_RBIT             : integer:=31;

--//���� C_HREG_IRQ_NUM - ������ ���������� ����������:
constant C_HIRQ_PCIE_DMA                      : integer:=0;
constant C_HIRQ_CFG_RX                        : integer:=1;
constant C_HIRQ_ETH_RX                        : integer:=2;
constant C_HIRQ_EDEV_RX                       : integer:=3;
constant C_HIRQ_PULT_RX                       : integer:=4;
constant C_HIRQ_VCH0                          : integer:=5;
constant C_HIRQ_VCH1                          : integer:=6;
constant C_HIRQ_VCH2                          : integer:=7;
constant C_HIRQ_VCH3                          : integer:=8;
constant C_HIRQ_VCH4                          : integer:=9;
constant C_HIRQ_VCH5                          : integer:=10;
constant C_HIRQ_VIZIR_RX                      : integer:=11;
constant C_HIRQ_BUP_RX                        : integer:=12;
constant C_HIRQ_PROM                          : integer:=13;
constant C_HIRQ_COUNT                         : integer:=C_HIRQ_PROM+1;
constant C_HIRQ_COUNT_MAX                     : integer:=pwr(2, (C_HREG_IRQ_NUM_M_WBIT-C_HREG_IRQ_NUM_L_WBIT+1));


--//Register C_HREG_MEM_ADR / Bit Map:
constant C_HREG_MEM_ADR_BANK_L_BIT            : integer:=31;--MEM_ADR_OFFSET[30..0]
constant C_HREG_MEM_ADR_BANK_M_BIT            : integer:=31;
constant C_HREG_MEM_ADR_LAST_BIT              : integer:=C_HREG_MEM_ADR_BANK_M_BIT;

--//Register C_HREG_MEM_CTRL / Bit Map:
constant C_HREG_MEM_CTRL_TRNWR_L_BIT          : integer:=0;
constant C_HREG_MEM_CTRL_TRNWR_M_BIT          : integer:=7;
constant C_HREG_MEM_CTRL_TRNRD_L_BIT          : integer:=8;
constant C_HREG_MEM_CTRL_TRNRD_M_BIT          : integer:=15;
constant C_HREG_MEM_CTRL_LAST_BIT             : integer:=C_HREG_MEM_CTRL_TRNRD_M_BIT;


--//Register C_HREG_PCIE / Bit Map:
--constant RESERV                             : integer:=5..0;
constant C_HREG_PCIE_NEG_LINK_L_RBIT          : integer:=6;
constant C_HREG_PCIE_NEG_LINK_M_RBIT          : integer:=11;
--constant RESERV                             : integer:=14...12;
constant C_HREG_PCIE_NEG_MAX_PAYLOAD_L_BIT    : integer:=15;
constant C_HREG_PCIE_NEG_MAX_PAYLOAD_M_BIT    : integer:=17;
constant C_HREG_PCIE_NEG_MAX_RD_REQ_L_BIT     : integer:=18;
constant C_HREG_PCIE_NEG_MAX_RD_REQ_M_BIT     : integer:=20;
--constant RESERV                             : integer:=27...21;
constant C_HREG_PCIE_SPEED_TESTING_BIT        : integer:=28;
constant C_HREG_PCIE_LAST_BIT                 : integer:=C_HREG_PCIE_SPEED_TESTING_BIT;


--//Register C_HREG_FUNC / Bit Map:
--//1/0 - ������������/�� ������������ � ������� FPGA
constant C_HREG_FUNC_MEM_BIT                  : integer:=0;
constant C_HREG_FUNC_TMR_BIT                  : integer:=1;
constant C_HREG_FUNC_VCTRL_BIT                : integer:=2;
constant C_HREG_FUNC_ETH_BIT                  : integer:=3;
constant C_HREG_FUNC_HDD_BIT                  : integer:=4;
constant C_HREG_FUNC_VRESEK21_BIT             : integer:=5;
constant C_HREG_FUNC_PROM_BIT                 : integer:=6;
constant C_HREG_FUNC_PULT_BIT                 : integer:=7;
constant C_HREG_FUNC_LAST_BIT                 : integer:=C_HREG_FUNC_PULT_BIT;


--//Register C_HREG_FUNCPRM / Bit Map:
constant C_HREG_FUNCPRM_MEMBANK_SIZE_L_BIT    : integer:=0;
constant C_HREG_FUNCPRM_MEMBANK_SIZE_M_BIT    : integer:=2;
constant C_HREG_FUNCPRM_VCTRL_VCH_COUNT_L_BIT : integer:=3;
constant C_HREG_FUNCPRM_VCTRL_VCH_COUNT_M_BIT : integer:=5;
constant C_HREG_FUNCPRM_VCTRL_MIR_BIT         : integer:=6;
constant C_HREG_FUNCPRM_LAST_BIT              : integer:=C_HREG_FUNCPRM_VCTRL_MIR_BIT;


--//���� ������ dsn_host.vhd /p_in_dev_option/ Bit Map:
constant C_HDEV_OPTIN_TXFIFO_PFULL_BIT        : integer:=0;
constant C_HDEV_OPTIN_RXFIFO_EMPTY_BIT        : integer:=1;
constant C_HDEV_OPTIN_MEMTRN_DONE_BIT         : integer:=2;
constant C_HDEV_OPTIN_VCTRL_FRMRK_L_BIT       : integer:=3;
constant C_HDEV_OPTIN_VCTRL_FRMRK_M_BIT       : integer:=34;
constant C_HDEV_OPTIN_VCTRL_FRSKIP_L_BIT      : integer:=35;
constant C_HDEV_OPTIN_VCTRL_FRSKIP_M_BIT      : integer:=42;
constant C_HDEV_OPTIN_TIME_L_BIT              : integer:=43;
constant C_HDEV_OPTIN_TIME_M_BIT              : integer:=74;
constant C_HDEV_OPTIN_LAST_BIT                : integer:=C_HDEV_OPTIN_TIME_M_BIT;

--//���� ������ dsn_host.vhd /p_out_dev_option/ Bit Map:
constant C_HDEV_OPTOUT_MEM_ADR_L_BIT          : integer:=0;
constant C_HDEV_OPTOUT_MEM_ADR_M_BIT          : integer:=31;
constant C_HDEV_OPTOUT_MEM_RQLEN_L_BIT        : integer:=32;
constant C_HDEV_OPTOUT_MEM_RQLEN_M_BIT        : integer:=49;--mem_rqlen: �������� � BYTE(max 128KB)
constant C_HDEV_OPTOUT_MEM_TRNWR_LEN_L_BIT    : integer:=50;
constant C_HDEV_OPTOUT_MEM_TRNWR_LEN_M_BIT    : integer:=57;--mem_trnwr: �������� � DWORD
constant C_HDEV_OPTOUT_MEM_TRNRD_LEN_L_BIT    : integer:=58;
constant C_HDEV_OPTOUT_MEM_TRNRD_LEN_M_BIT    : integer:=65;--mem_trnrd: �������� � DWORD
constant C_HDEV_OPTOUT_TIME_L_BIT             : integer:=66;
constant C_HDEV_OPTOUT_TIME_M_BIT             : integer:=97;
constant C_HDEV_OPTOUT_TIME_SET_BIT           : integer:=98;
constant C_HDEV_OPTOUT_LAST_BIT               : integer:=C_HDEV_OPTOUT_TIME_SET_BIT;



--//--------------------------------------------------------------
--//������ ���������������� (cfgdev.vhd)
--//--------------------------------------------------------------
--//������ ��������� ��������� ����� ������ cfgdev.vhd
--//Device Address map:
constant C_CFGDEV_SWT                         : integer:=16#00#;
constant C_CFGDEV_ETH                         : integer:=16#01#;
constant C_CFGDEV_VCTRL                       : integer:=16#02#;
constant C_CFGDEV_TMR                         : integer:=16#03#;
--constant RESERV                               : integer:=16#04#;
constant C_CFGDEV_HDD                         : integer:=16#05#;
constant C_CFGDEV_TESTING                     : integer:=16#06#;
constant C_CFGDEV_COUNT                       : integer:=C_CFGDEV_TESTING + 1;
constant C_CFGDEV_COUNT_MAX                   : integer:=256;--������������ ����������� C_CFGPKT_DADR_M/L_BIT � cfgdev_pkg.vhd



--//--------------------------------------------------------------
--//�������� ������ dsn_timer.vhd
--//--------------------------------------------------------------
constant C_TMR_REG_CTRL                       : integer:=16#000#;
constant C_TMR_REG_CMP_L                      : integer:=16#001#;
constant C_TMR_REG_CMP_M                      : integer:=16#002#;


--//Register C_TMR_REG_CTRL / Bit Map:
constant C_TMR_REG_CTRL_NUM_L_BIT             : integer:=0;--����� �������
constant C_TMR_REG_CTRL_NUM_M_BIT             : integer:=3;
constant C_TMR_REG_CTRL_EN_BIT                : integer:=14;
constant C_TMR_REG_CTRL_DIS_BIT               : integer:=15;
--constant C_TMR_REG_CTRL_STATUS_EN_L_RBIT      : integer:=0;--������ ��� ������ ���. C_TMR_REG_CTRL
--constant C_TMR_REG_CTRL_STATUS_EN_M_RBIT      : integer:=xxx;
constant C_TMR_REG_CTRL_LAST_BIT              : integer:=C_TMR_REG_CTRL_DIS_BIT;


--//���������� ���-�� �������� � dsn_timer.vhd
constant C_TMR_COUNT                          : integer:=6;
constant C_TMR_COUNT_MAX                      : integer:=pwr(2, (C_TMR_REG_CTRL_NUM_M_BIT-C_TMR_REG_CTRL_NUM_L_BIT+1));

constant C_TMR_ETH                            : integer:=0;
constant C_TMR_EDEV                           : integer:=1;
constant C_TMR_PULT                           : integer:=2;
constant C_TMR_BUP                            : integer:=3;
constant C_TMR_VIZIR                          : integer:=4;


--//--------------------------------------------------------------
--//�������� ������ dsn_switch.vhd
--//--------------------------------------------------------------
constant C_SWT_REG_CTRL                       : integer:=16#07#;
constant C_SWT_REG_FRR_ETHG_HOST              : integer:=16#08#;
constant C_SWT_REG_FRR_ETHG_VCTRL             : integer:=16#10#;
constant C_SWT_REG_FRR_ETHG_HDD               : integer:=16#18#;


--//Register C_SWT_REG_CTRL / Bit Map:
constant C_SWT_REG_CTRL_RST_ETH_BUFS_BIT      : integer:=0;
constant C_SWT_REG_CTRL_RST_VCTRL_BUFS_BIT    : integer:=1;
constant C_SWT_REG_CTRL_TSTDSN_2_ETHTXBUF_BIT : integer:=2;
constant C_SWT_REG_CTRL_LAST_BIT              : integer:=C_SWT_REG_CTRL_TSTDSN_2_ETHTXBUF_BIT;


--//��� ���-�� ������ �������������:
constant C_SWT_FRR_COUNT_MAX                  : integer:=8;

--//
constant C_SWT_ETH_HOST_FRR_COUNT             : integer:=3;--���-�� ������ ������������ ������� ETH-HOST
constant C_SWT_ETH_VCTRL_FRR_COUNT            : integer:=C_PCFG_VCTRL_VCH_COUNT;--���-�� ������ ������������ ������� ETH-VCTRL
constant C_SWT_ETH_HDD_FRR_COUNT              : integer:=3;--//���-�� ������ ������������ ������� ETH-HDD

Type TEthFRRGet is array (0 to C_SWT_FRR_COUNT_MAX-1) of integer;
----------------------------------------------------------------------------------------
--//C_SWT_ETH_xxx_FRR_COUNT - ��������:          | 1 | 2 | 3 | 4 | 5 | 6 | 7 | 8 |
----------------------------------------------------------------------------------------
constant C_SWT_GET_FMASK_REG_COUNT : TEthFRRGet:=( 1,  1,  2,  2,  3,  3,  4,  4 );
Type TEthFRR is array (0 to C_SWT_FRR_COUNT_MAX-1) of std_logic_vector(7 downto 0);
--����� ���������� (7...0), ���
-- 3..0 - ��� ������
-- 7..4 - ������ ������



--//--------------------------------------------------------------
--//�������� ������ dsn_eth.vhd
--//--------------------------------------------------------------
constant C_ETH_REG_CTRL                       : integer:=16#000#;
constant C_ETH_REG_MAC_PATRN0                 : integer:=16#001#;--DST MAC
constant C_ETH_REG_MAC_PATRN1                 : integer:=16#002#;
constant C_ETH_REG_MAC_PATRN2                 : integer:=16#003#;
constant C_ETH_REG_MAC_PATRN3                 : integer:=16#004#;--SRC MAC
constant C_ETH_REG_MAC_PATRN4                 : integer:=16#005#;
constant C_ETH_REG_MAC_PATRN5                 : integer:=16#006#;
constant C_ETH_REG_IP_PATRN0                  : integer:=16#007#;--DST IP
constant C_ETH_REG_IP_PATRN1                  : integer:=16#008#;
constant C_ETH_REG_IP_PATRN2                  : integer:=16#009#;--SRC IP
constant C_ETH_REG_IP_PATRN3                  : integer:=16#00A#;
constant C_ETH_REG_PORT_PATRN0                : integer:=16#00B#;--DST PORT
constant C_ETH_REG_PORT_PATRN1                : integer:=16#00C#;--SRC PORT


--//--------------------------------------------------------------
--//�������� ������ dsn_video_ctrl.vhd
--//--------------------------------------------------------------
constant C_VCTRL_REG_CTRL                     : integer:=16#000#;
constant C_VCTRL_REG_DATA_L                   : integer:=16#001#;
constant C_VCTRL_REG_DATA_M                   : integer:=16#002#;
constant C_VCTRL_REG_MEM_CTRL                 : integer:=16#003#;--(15..8)(7..0) - trn_mem_rd;trn_mem_wr
constant C_VCTRL_REG_TST0                     : integer:=16#004#;


--//Register C_VCTRL_REG_CTRL / Bit Map:
constant C_VCTRL_REG_CTRL_VCH_L_BIT           : integer:=0; --����� ����� ������
constant C_VCTRL_REG_CTRL_VCH_M_BIT           : integer:=3;
constant C_VCTRL_REG_CTRL_PRM_L_BIT           : integer:=4; --����� ��������
constant C_VCTRL_REG_CTRL_PRM_M_BIT           : integer:=6;
constant C_VCTRL_REG_CTRL_SET_BIT             : integer:=7;
constant C_VCTRL_REG_CTRL_SET_IDLE_BIT        : integer:=8;
constant C_VCTRL_REG_CTRL_RAMCOE_ADR_BIT      : integer:=9;
constant C_VCTRL_REG_CTRL_RAMCOE_DATA_BIT     : integer:=10;
constant C_VCTRL_REG_CTRL_RAMCOE_L_BIT        : integer:=11;--����� RAMCOE
constant C_VCTRL_REG_CTRL_RAMCOE_M_BIT        : integer:=14;
constant C_VCTRL_REG_CTRL_LAST_BIT            : integer:=C_VCTRL_REG_CTRL_RAMCOE_M_BIT;

--//������� ��� ���� VCTRL_REG_CTRL_RAMCOENUM:
constant C_VCTRL_RAMCOE_SCALE                 : integer:=0;
constant C_VCTRL_RAMCOE_PCOLR                 : integer:=1;
constant C_VCTRL_RAMCOE_PCOLG                 : integer:=2;
constant C_VCTRL_RAMCOE_PCOLB                 : integer:=3;
constant C_VCTRL_RAMCOE_GAMMA_GRAY            : integer:=4;
constant C_VCTRL_RAMCOE_GAMMA_COLR            : integer:=5;
constant C_VCTRL_RAMCOE_GAMMA_COLG            : integer:=6;
constant C_VCTRL_RAMCOE_GAMMA_COLB            : integer:=7;

--//������� ��� ���� VCTRL_REG_CTRL_PRMNUM:
constant C_VCTRL_PRM_MEM_ADR_WR               : integer:=0;--������� ����� ������ ������ �����
constant C_VCTRL_PRM_MEM_ADR_RD               : integer:=1;--������� ����� ������ ������ �����
constant C_VCTRL_PRM_FR_ZONE_SKIP             : integer:=2;
constant C_VCTRL_PRM_FR_ZONE_ACTIVE           : integer:=3;
constant C_VCTRL_PRM_FR_OPTIONS               : integer:=4;
--//��� ���-�� ������� ��������� ����������:
constant C_VCTRL_PRM_COUNT_MAX                : integer:=pwr(2, (C_VCTRL_REG_CTRL_PRM_M_BIT-C_VCTRL_REG_CTRL_PRM_L_BIT+1));


--//Register VCTRL_REG_MEM_ADDR / Bit Map:
constant C_VCTRL_REG_MEM_ADR_BANK_L_BIT       : integer:=C_HREG_MEM_ADR_BANK_L_BIT;
constant C_VCTRL_REG_MEM_ADR_BANK_M_BIT       : integer:=C_HREG_MEM_ADR_BANK_M_BIT;
constant C_VCTRL_REG_MEM_LAST_BIT             : integer:=C_VCTRL_REG_MEM_ADR_BANK_M_BIT;

--//Memory map for video: (max frame size: 2048x2048)
--//                                          : integer:=0; --������� ����������(VLINE_LSB-1...0)
constant C_VCTRL_MEM_VLINE_L_BIT              : integer:=C_PCFG_VCTRL_MEM_VLINE_L_BIT;--������ ���������� (MSB...LSB)
constant C_VCTRL_MEM_VLINE_M_BIT              : integer:=C_PCFG_VCTRL_MEM_VLINE_M_BIT;
constant C_VCTRL_MEM_VFR_L_BIT                : integer:=C_PCFG_VCTRL_MEM_VFR_L_BIT  ;--����� ����� (MSB...LSB) - �����������
constant C_VCTRL_MEM_VFR_M_BIT                : integer:=C_PCFG_VCTRL_MEM_VFR_M_BIT  ;
constant C_VCTRL_MEM_VCH_L_BIT                : integer:=C_PCFG_VCTRL_MEM_VCH_L_BIT  ;--����� ����� ������ (MSB...LSB)
constant C_VCTRL_MEM_VCH_M_BIT                : integer:=C_PCFG_VCTRL_MEM_VCH_M_BIT  ;

--//��� ���-�� ����� �������:
constant C_VCTRL_VCH_COUNT                    : integer:=C_PCFG_VCTRL_VCH_COUNT;
constant C_VCTRL_VCH_COUNT_MAX                : integer:=pwr(2, (C_VCTRL_MEM_VCH_M_BIT-C_VCTRL_MEM_VCH_L_BIT+1));


--//Register C_VCTRL_REG_TST0 / Bit Map:
constant C_VCTRL_REG_TST0_DBG_TBUFRD_BIT      : integer:=0;--������� ������ �������� - ����������� ����������� RAM/TRACK/TBUF
constant C_VCTRL_REG_TST0_DBG_EBUFRD_BIT      : integer:=1;--������� ������ �������� - ����������� ����������� RAM/TRACK/EBUF
constant C_VCTRL_REG_TST0_DBG_SOBEL_BIT       : integer:=2;--1/0 - ������� ������ ������ ������ Grad/Video
constant C_VCTRL_REG_TST0_DBG_ROTRIGHT_BIT    : integer:=3;--������� �� 90 ������
constant C_VCTRL_REG_TST0_DBG_ROTLEFT_BIT     : integer:=4;--������� �� 90 �����
constant C_VCTRL_REG_TST0_DBG_DIS_DEMCOLOR_BIT: integer:=5;--1/0 - ��������� ������ ������ vcoldemosaic_main.vhd
constant C_VCTRL_REG_TST0_DBG_DCOUNT_BIT      : integer:=6;--1 - ������ ������ ������ ����������� �������
constant C_VCTRL_REG_TST0_DBG_PICTURE_BIT     : integer:=7;--�������� ������ ����� � ��� + �������� ������������� �������� vbuf,
                                                           --��� ���(7)=1 - vbuf=0
constant C_VCTRL_REG_TST0_SKIPFR_CNT_CLR_BIT  : integer:=8;--��� 1 - ���������� ����� ��������� ���������� ������ tst_vfrskip,
                                                           --��� 0 - ���
--constant RESERV                               : integer:=9;
constant C_VCTRL_REG_TST0_DBG_RDHOLD_BIT      : integer:=10;--�������� ������� ����������� ������� ������
constant C_VCTRL_REG_TST0_DBG_TRCHOLD_BIT     : integer:=11;--�������� ������� ����������� ������� ��������
constant C_VCTRL_REG_TST0_LAST_BIT            : integer:=C_VCTRL_REG_TST0_DBG_TRCHOLD_BIT;



end prj_def;


package body prj_def is

end prj_def;

