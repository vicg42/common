-------------------------------------------------------------------------
-- Company     : Telemix
-- Engineer    : Golovachenko Victor
--
-- Create Date : 10/26/2007
-- Module Name :
--
-- Description :
--
-- Revision:
-- Revision 0.01 - File Created
--
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
-- need conversion function to convert reals/integers to std logic vectors
use ieee.std_logic_arith.conv_std_logic_vector;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


package test_im_pkg is


type TBmp_FileHeader is record
bfType      : std_logic_vector(15 downto 0);--WORD
bfSize      : std_logic_vector(31 downto 0);--DWORD
bfReserved1 : std_logic_vector(15 downto 0);--WORD
bfReserved2 : std_logic_vector(15 downto 0);--WORD
bfOffBits   : std_logic_vector(31 downto 0);--DWORD
end record;

type TBmp_InfoHeader is record
biSize         : std_logic_vector(31 downto 0);--DWORD
biWidth        : std_logic_vector(63 downto 0);--LONG
biHeight       : std_logic_vector(63 downto 0);--LONG
biPlanes       : std_logic_vector(15 downto 0);--WORD
biBitCount     : std_logic_vector(15 downto 0);--WORD
biCompression  : std_logic_vector(31 downto 0);--DWORD
biSizeImage    : std_logic_vector(31 downto 0);--DWORD
biXPelsPerMeter: std_logic_vector(63 downto 0);--LONG
biYPelsPerMeter: std_logic_vector(63 downto 0);--LONG
biClrUsed      : std_logic_vector(31 downto 0);--DWORD
biClrImportant : std_logic_vector(31 downto 0);--DWORD
end record;

type TBmp_Info is record
fh : TBmp_FileHeader;
ih : TBmp_InfoHeader;
end record;


--//�������� �������� - tst.png (24x16)
type TImageTst  is array (0 to (8*17)-1) of std_logic_vector (31 downto 0);
constant IMAGE_TST00 : TImageTst:=(
--//Y0
(CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#017#, 8)&CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#178#, 8)&CONV_STD_LOGIC_VECTOR(10#163#, 8)&CONV_STD_LOGIC_VECTOR(10#096#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#117#, 8)&CONV_STD_LOGIC_VECTOR(10#157#, 8)&CONV_STD_LOGIC_VECTOR(10#160#, 8)&CONV_STD_LOGIC_VECTOR(10#161#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y1
(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#053#, 8)&CONV_STD_LOGIC_VECTOR(10#086#, 8)&CONV_STD_LOGIC_VECTOR(10#047#, 8)&CONV_STD_LOGIC_VECTOR(10#017#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#036#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#172#, 8)&CONV_STD_LOGIC_VECTOR(10#174#, 8)&CONV_STD_LOGIC_VECTOR(10#119#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#107#, 8)&CONV_STD_LOGIC_VECTOR(10#152#, 8)&CONV_STD_LOGIC_VECTOR(10#157#, 8)&CONV_STD_LOGIC_VECTOR(10#155#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y2
(CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#135#, 8)&CONV_STD_LOGIC_VECTOR(10#077#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#179#, 8)&CONV_STD_LOGIC_VECTOR(10#234#, 8)&CONV_STD_LOGIC_VECTOR(10#190#, 8)&CONV_STD_LOGIC_VECTOR(10#152#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)&CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#068#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#179#, 8)&CONV_STD_LOGIC_VECTOR(10#195#, 8)&CONV_STD_LOGIC_VECTOR(10#159#, 8)&CONV_STD_LOGIC_VECTOR(10#045#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#076#, 8)&CONV_STD_LOGIC_VECTOR(10#132#, 8)&CONV_STD_LOGIC_VECTOR(10#154#, 8)&CONV_STD_LOGIC_VECTOR(10#161#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y3
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)&CONV_STD_LOGIC_VECTOR(10#016#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#227#, 8)&CONV_STD_LOGIC_VECTOR(10#107#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#032#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#242#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#243#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#009#, 8)&CONV_STD_LOGIC_VECTOR(10#007#, 8)&CONV_STD_LOGIC_VECTOR(10#063#, 8)&CONV_STD_LOGIC_VECTOR(10#169#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#219#, 8)&CONV_STD_LOGIC_VECTOR(10#235#, 8)&CONV_STD_LOGIC_VECTOR(10#211#, 8)&CONV_STD_LOGIC_VECTOR(10#087#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#064#, 8)&CONV_STD_LOGIC_VECTOR(10#136#, 8)&CONV_STD_LOGIC_VECTOR(10#187#, 8)&CONV_STD_LOGIC_VECTOR(10#207#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y4
(CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#191#, 8)&CONV_STD_LOGIC_VECTOR(10#074#, 8)&CONV_STD_LOGIC_VECTOR(10#049#, 8)&CONV_STD_LOGIC_VECTOR(10#058#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#247#, 8)&CONV_STD_LOGIC_VECTOR(10#230#, 8)&CONV_STD_LOGIC_VECTOR(10#248#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#053#, 8)&CONV_STD_LOGIC_VECTOR(10#164#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#247#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)&CONV_STD_LOGIC_VECTOR(10#119#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#067#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y5
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#097#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#043#, 8)&CONV_STD_LOGIC_VECTOR(10#053#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#243#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#217#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#074#, 8)&CONV_STD_LOGIC_VECTOR(10#143#, 8)&CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#245#, 8)&CONV_STD_LOGIC_VECTOR(10#248#, 8)&CONV_STD_LOGIC_VECTOR(10#245#, 8)&CONV_STD_LOGIC_VECTOR(10#148#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#058#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#244#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y6
(CONV_STD_LOGIC_VECTOR(10#013#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#047#, 8)&CONV_STD_LOGIC_VECTOR(10#042#, 8)&CONV_STD_LOGIC_VECTOR(10#077#, 8)&CONV_STD_LOGIC_VECTOR(10#055#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#238#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)&CONV_STD_LOGIC_VECTOR(10#157#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#162#, 8)&CONV_STD_LOGIC_VECTOR(10#214#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#249#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)&CONV_STD_LOGIC_VECTOR(10#253#, 8)&CONV_STD_LOGIC_VECTOR(10#200#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#050#, 8)&CONV_STD_LOGIC_VECTOR(10#139#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#253#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y7
(CONV_STD_LOGIC_VECTOR(10#028#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)&CONV_STD_LOGIC_VECTOR(10#025#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#065#, 8)&CONV_STD_LOGIC_VECTOR(10#127#, 8)&CONV_STD_LOGIC_VECTOR(10#172#, 8)&CONV_STD_LOGIC_VECTOR(10#106#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#249#, 8)&CONV_STD_LOGIC_VECTOR(10#251#, 8)&CONV_STD_LOGIC_VECTOR(10#205#, 8)&CONV_STD_LOGIC_VECTOR(10#091#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#221#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)&CONV_STD_LOGIC_VECTOR(10#247#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#239#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#048#, 8)&CONV_STD_LOGIC_VECTOR(10#120#, 8)&CONV_STD_LOGIC_VECTOR(10#216#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y8
(CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#009#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#013#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#159#, 8)&CONV_STD_LOGIC_VECTOR(10#199#, 8)&CONV_STD_LOGIC_VECTOR(10#198#, 8)&CONV_STD_LOGIC_VECTOR(10#107#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#226#, 8)&CONV_STD_LOGIC_VECTOR(10#143#, 8)&CONV_STD_LOGIC_VECTOR(10#105#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#228#, 8)&CONV_STD_LOGIC_VECTOR(10#237#, 8)&CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#247#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#239#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)&CONV_STD_LOGIC_VECTOR(10#248#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#125#, 8)&CONV_STD_LOGIC_VECTOR(10#144#, 8)&CONV_STD_LOGIC_VECTOR(10#237#, 8)&CONV_STD_LOGIC_VECTOR(10#252#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y9
(CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#032#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#175#, 8)&CONV_STD_LOGIC_VECTOR(10#165#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#091#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#219#, 8)&CONV_STD_LOGIC_VECTOR(10#158#, 8)&CONV_STD_LOGIC_VECTOR(10#127#, 8)&CONV_STD_LOGIC_VECTOR(10#154#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#220#, 8)&CONV_STD_LOGIC_VECTOR(10#235#, 8)&CONV_STD_LOGIC_VECTOR(10#254#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#252#, 8)&CONV_STD_LOGIC_VECTOR(10#253#, 8)&CONV_STD_LOGIC_VECTOR(10#250#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#145#, 8)&CONV_STD_LOGIC_VECTOR(10#121#, 8)&CONV_STD_LOGIC_VECTOR(10#211#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y10
(CONV_STD_LOGIC_VECTOR(10#015#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#034#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#181#, 8)&CONV_STD_LOGIC_VECTOR(10#184#, 8)&CONV_STD_LOGIC_VECTOR(10#187#, 8)&CONV_STD_LOGIC_VECTOR(10#100#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#183#, 8)&CONV_STD_LOGIC_VECTOR(10#136#, 8)&CONV_STD_LOGIC_VECTOR(10#144#, 8)&CONV_STD_LOGIC_VECTOR(10#183#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#212#, 8)&CONV_STD_LOGIC_VECTOR(10#233#, 8)&CONV_STD_LOGIC_VECTOR(10#249#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#254#, 8)&CONV_STD_LOGIC_VECTOR(10#242#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#102#, 8)&CONV_STD_LOGIC_VECTOR(10#084#, 8)&CONV_STD_LOGIC_VECTOR(10#175#, 8)&CONV_STD_LOGIC_VECTOR(10#246#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y11
(CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#038#, 8)&CONV_STD_LOGIC_VECTOR(10#019#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#195#, 8)&CONV_STD_LOGIC_VECTOR(10#228#, 8)&CONV_STD_LOGIC_VECTOR(10#218#, 8)&CONV_STD_LOGIC_VECTOR(10#090#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#202#, 8)&CONV_STD_LOGIC_VECTOR(10#204#, 8)&CONV_STD_LOGIC_VECTOR(10#217#, 8)&CONV_STD_LOGIC_VECTOR(10#215#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#220#, 8)&CONV_STD_LOGIC_VECTOR(10#236#, 8)&CONV_STD_LOGIC_VECTOR(10#232#, 8)&CONV_STD_LOGIC_VECTOR(10#218#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#217#, 8)&CONV_STD_LOGIC_VECTOR(10#216#, 8)&CONV_STD_LOGIC_VECTOR(10#207#, 8)&CONV_STD_LOGIC_VECTOR(10#226#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#131#, 8)&CONV_STD_LOGIC_VECTOR(10#131#, 8)&CONV_STD_LOGIC_VECTOR(10#168#, 8)&CONV_STD_LOGIC_VECTOR(10#198#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y12
(CONV_STD_LOGIC_VECTOR(10#010#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#040#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#140#, 8)&CONV_STD_LOGIC_VECTOR(10#152#, 8)&CONV_STD_LOGIC_VECTOR(10#130#, 8)&CONV_STD_LOGIC_VECTOR(10#039#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#185#, 8)&CONV_STD_LOGIC_VECTOR(10#183#, 8)&CONV_STD_LOGIC_VECTOR(10#174#, 8)&CONV_STD_LOGIC_VECTOR(10#148#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#202#, 8)&CONV_STD_LOGIC_VECTOR(10#206#, 8)&CONV_STD_LOGIC_VECTOR(10#192#, 8)&CONV_STD_LOGIC_VECTOR(10#182#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#172#, 8)&CONV_STD_LOGIC_VECTOR(10#165#, 8)&CONV_STD_LOGIC_VECTOR(10#150#, 8)&CONV_STD_LOGIC_VECTOR(10#175#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#206#, 8)&CONV_STD_LOGIC_VECTOR(10#206#, 8)&CONV_STD_LOGIC_VECTOR(10#187#, 8)&CONV_STD_LOGIC_VECTOR(10#167#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y13
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#034#, 8)&CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#024#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#046#, 8)&CONV_STD_LOGIC_VECTOR(10#036#, 8)&CONV_STD_LOGIC_VECTOR(10#033#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#088#, 8)&CONV_STD_LOGIC_VECTOR(10#067#, 8)&CONV_STD_LOGIC_VECTOR(10#055#, 8)&CONV_STD_LOGIC_VECTOR(10#041#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#146#, 8)&CONV_STD_LOGIC_VECTOR(10#128#, 8)&CONV_STD_LOGIC_VECTOR(10#108#, 8)&CONV_STD_LOGIC_VECTOR(10#094#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#144#, 8)&CONV_STD_LOGIC_VECTOR(10#156#, 8)&CONV_STD_LOGIC_VECTOR(10#143#, 8)&CONV_STD_LOGIC_VECTOR(10#135#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#216#, 8)&CONV_STD_LOGIC_VECTOR(10#224#, 8)&CONV_STD_LOGIC_VECTOR(10#193#, 8)&CONV_STD_LOGIC_VECTOR(10#153#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y14
(CONV_STD_LOGIC_VECTOR(10#026#, 8)&CONV_STD_LOGIC_VECTOR(10#020#, 8)&CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#030#, 8)&CONV_STD_LOGIC_VECTOR(10#021#, 8)&CONV_STD_LOGIC_VECTOR(10#027#, 8)&CONV_STD_LOGIC_VECTOR(10#023#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#022#, 8)&CONV_STD_LOGIC_VECTOR(10#008#, 8)&CONV_STD_LOGIC_VECTOR(10#012#, 8)&CONV_STD_LOGIC_VECTOR(10#018#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#091#, 8)&CONV_STD_LOGIC_VECTOR(10#050#, 8)&CONV_STD_LOGIC_VECTOR(10#035#, 8)&CONV_STD_LOGIC_VECTOR(10#028#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#128#, 8)&CONV_STD_LOGIC_VECTOR(10#180#, 8)&CONV_STD_LOGIC_VECTOR(10#179#, 8)&CONV_STD_LOGIC_VECTOR(10#151#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#157#, 8)&CONV_STD_LOGIC_VECTOR(10#166#, 8)&CONV_STD_LOGIC_VECTOR(10#129#, 8)&CONV_STD_LOGIC_VECTOR(10#104#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//28..31

--//Y15
(CONV_STD_LOGIC_VECTOR(10#029#, 8)&CONV_STD_LOGIC_VECTOR(10#014#, 8)&CONV_STD_LOGIC_VECTOR(10#011#, 8)&CONV_STD_LOGIC_VECTOR(10#005#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#041#, 8)&CONV_STD_LOGIC_VECTOR(10#039#, 8)&CONV_STD_LOGIC_VECTOR(10#038#, 8)&CONV_STD_LOGIC_VECTOR(10#029#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#075#, 8)&CONV_STD_LOGIC_VECTOR(10#047#, 8)&CONV_STD_LOGIC_VECTOR(10#040#, 8)&CONV_STD_LOGIC_VECTOR(10#041#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#113#, 8)&CONV_STD_LOGIC_VECTOR(10#064#, 8)&CONV_STD_LOGIC_VECTOR(10#071#, 8)&CONV_STD_LOGIC_VECTOR(10#084#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#189#, 8)&CONV_STD_LOGIC_VECTOR(10#255#, 8)&CONV_STD_LOGIC_VECTOR(10#240#, 8)&CONV_STD_LOGIC_VECTOR(10#206#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#105#, 8)&CONV_STD_LOGIC_VECTOR(10#114#, 8)&CONV_STD_LOGIC_VECTOR(10#082#, 8)&CONV_STD_LOGIC_VECTOR(10#104#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)),  --//28..31


--//Y16
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//0..3
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//4..7
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//8..11
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//12..15
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//16..19
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//20..23
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)), --//24..27
(CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8)&CONV_STD_LOGIC_VECTOR(10#000#, 8))  --//28..31

);

end test_im_pkg;

package body test_im_pkg is


end package body test_im_pkg;

