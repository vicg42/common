-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 20.01.2013 15:47:02
-- Module Name : clocks
--
-- ����������/�������� :
--
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.clocks_pkg.all;
use work.prj_cfg.all;

entity clocks is
port(
p_out_rst  : out   std_logic;
p_out_gclk : out   std_logic_vector(7 downto 0);

p_in_clkopt: in    std_logic_vector(3 downto 0);
p_in_clk   : in    TRefClkPinIN
);
end;

architecture synth of clocks is

signal i_pll_clkin   : std_logic;
signal g_pll_clkin   : std_logic;
signal i_pll_rst_cnt : std_logic_vector(4 downto 0) := "11111";
signal i_pll_rst     : std_logic := '1';
signal i_clk_fb      : std_logic_vector(2 downto 0);
signal g_clk_fb      : std_logic_vector(2 downto 0);
signal i_pll_locked  : std_logic_vector(2 downto 0);
signal i_clk_out     : std_logic_vector(7 downto 0);
signal g_clk         : std_logic_vector(7 downto 0);

begin

m_buf : IBUFDS port map(I  => p_in_clk.clk_p, IB => p_in_clk.clk_n, O => i_pll_clkin);--200MHz
bufg_pll_clkin : BUFG port map(I  => i_pll_clkin, O  => g_pll_clkin);

process(g_pll_clkin)
begin
  if rising_edge(g_pll_clkin) then
    if i_pll_rst_cnt = "00000" then
      i_pll_rst <= '0';
    else
      i_pll_rst <= '1';
      i_pll_rst_cnt <= i_pll_rst_cnt-1;
    end if;
  end if;
end process;

-- Generate asynchronous reset
p_out_rst <= not(OR_reduce(i_pll_locked));

p_out_gclk(0) <= g_pll_clkin;
bufg_clk1: BUFG port map(I => i_clk_out(1), O => p_out_gclk(1)); --300MHz
bufg_clk2: BUFG port map(I => i_clk_out(0), O => g_clk(0)); p_out_gclk(2) <= g_clk(0); --100MHz
m_buf_pciexp : IBUFDS port map(I  => p_in_clk.pciexp_clk_p, IB => p_in_clk.pciexp_clk_n, O => p_out_gclk(3));
bufg_clk4: BUFG port map(I => i_clk_out(4), O => g_clk(4)); p_out_gclk(4) <= g_clk(4); --125MHz
bufg_clk5: BUFG port map(I => i_clk_out(5), O => p_out_gclk(5));--65,625MHz
p_out_gclk(6) <= g_pll_clkin;--200MHz   --bufg_clk6: BUFG port map(I => i_clk_out(2), O => p_out_gclk(6));--450 MHz
p_out_gclk(7 downto 7)<=(others=>'0');

-- Reference clock PLL (CLKFBOUT range 400 MHz to 1000 MHz)
-- CLKFBOUT = (CLKIN1/DIVCLK_DIVIDE) * CLKFBOUT_MULT
-- CLKOUTn  = (CLKIN1/DIVCLK_DIVIDE) * CLKFBOUT_MULT/CLKOUTn_DIVIDE
-- CLKFBOUT = (200 MHz/2) * 9.000       = 900 MHz
-- CLKOUT0  = (200 MHz/2) * 9.000/9     = 100 MHz
-- CLKOUT1  = (200 MHz/2) * 9.000/3     = 300 MHz (mem_clk)
-- CLKOUT2  = (200 MHz/2) * 9.000/2     = 450 MHz

m_pll0 : PLL_BASE
generic map(
CLKIN_PERIOD   => 5.00,  --200MHz
DIVCLK_DIVIDE  => 2,     --integer : 1 to 52
CLKFBOUT_MULT  => 9,     --integer : 1 to 64
CLKOUT0_DIVIDE => 9,     --integer : 1 to 128
CLKOUT1_DIVIDE => 3,     --integer : 1 to 128
CLKOUT2_DIVIDE => 2,     --integer : 1 to 128
CLKOUT3_DIVIDE => 1,     --integer : 1 to 128
CLKOUT0_PHASE  => 0.000,
CLKOUT1_PHASE  => 0.000,
CLKOUT2_PHASE  => 0.000,
CLKOUT3_PHASE  => 0.000
)
port map(
CLKFBOUT => i_clk_fb(0),
CLKOUT0  => i_clk_out(0),
CLKOUT1  => i_clk_out(1),
CLKOUT2  => i_clk_out(2),
CLKOUT3  => open,
CLKOUT4  => open,
CLKOUT5  => open,
LOCKED   => i_pll_locked(0),
CLKFBIN  => g_clk_fb(0),
CLKIN    => i_pll_clkin,
RST      => i_pll_rst
);
-- MMCM feedback (not using BUFG, because we don't care about phase compensation)
g_clk_fb(0) <= i_clk_fb(0);


-- Reference clock PLL (CLKFBOUT range 400 MHz to 1000 MHz)
-- CLKFBOUT = (CLKIN1/DIVCLK_DIVIDE) * CLKFBOUT_MULT
-- CLKOUTn  = (CLKIN1/DIVCLK_DIVIDE) * CLKFBOUT_MULT/CLKOUTn_DIVIDE
-- CLKFBOUT = (100 MHz/1) * 5.000       = 500 MHz
-- CLKOUT0  = (100 MHz/1) * 5.000/4     = 125 MHz

m_pll1 : PLL_BASE
generic map(
CLKIN_PERIOD   => 10.00, --100MHz
DIVCLK_DIVIDE  => 1,     --integer : 1 to 52
CLKFBOUT_MULT  => 5,     --integer : 1 to 64
CLKOUT0_DIVIDE => 4,     --integer : 1 to 128
CLKOUT1_DIVIDE => 1,     --integer : 1 to 128
CLKOUT2_DIVIDE => 1,     --integer : 1 to 128
CLKOUT3_DIVIDE => 1,     --integer : 1 to 128
CLKOUT0_PHASE  => 0.000,
CLKOUT1_PHASE  => 0.000,
CLKOUT2_PHASE  => 0.000,
CLKOUT3_PHASE  => 0.000
)
port map(
CLKFBOUT => i_clk_fb(1),
CLKOUT0  => i_clk_out(4),
CLKOUT1  => open,
CLKOUT2  => open,
CLKOUT3  => open,
CLKOUT4  => open,
CLKOUT5  => open,
LOCKED   => i_pll_locked(1),
CLKFBIN  => g_clk_fb(1),
CLKIN    => g_clk(0),--i_clk_out(0),
RST      => i_pll_rst
);
-- MMCM feedback (not using BUFG, because we don't care about phase compensation)
g_clk_fb(1) <= i_clk_fb(1);


-- Reference clock PLL (CLKFBOUT range 400 MHz to 1000 MHz)
-- CLKFBOUT = (CLKIN1/DIVCLK_DIVIDE) * CLKFBOUT_MULT
-- CLKOUTn  = (CLKIN1/DIVCLK_DIVIDE) * CLKFBOUT_MULT/CLKOUTn_DIVIDE
-- CLKFBOUT = (125 MHz/4) * 21.000      = 656,25 MHz
-- CLKOUT0  = (125 MHz/4) * 21.000/10   = 65,625 MHz

m_pll2 : PLL_BASE
generic map(
CLKIN_PERIOD   => 8.00,  --125MHz
DIVCLK_DIVIDE  => 4,     --integer : 1 to 52
CLKFBOUT_MULT  => 21,    --integer : 1 to 64
CLKOUT0_DIVIDE => 10,    --integer : 1 to 128
CLKOUT1_DIVIDE => 1,     --integer : 1 to 128
CLKOUT2_DIVIDE => 1,     --integer : 1 to 128
CLKOUT3_DIVIDE => 1,     --integer : 1 to 128
CLKOUT0_PHASE  => 0.000,
CLKOUT1_PHASE  => 0.000,
CLKOUT2_PHASE  => 0.000,
CLKOUT3_PHASE  => 0.000
)
port map(
CLKFBOUT => i_clk_fb(2),
CLKOUT0  => i_clk_out(5),
CLKOUT1  => open,
CLKOUT2  => open,
CLKOUT3  => open,
CLKOUT4  => open,
CLKOUT5  => open,
LOCKED   => i_pll_locked(2),
CLKFBIN  => g_clk_fb(2),
CLKIN    => g_clk(4),
RST      => i_pll_rst
);
-- MMCM feedback (not using BUFG, because we don't care about phase compensation)
g_clk_fb(2) <= i_clk_fb(2);

end;