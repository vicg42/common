`timescale 1ns / 1ps
module cubic_table #(
    parameter PIXEL_STEP = 4096,
    parameter COE_WIDTH = 10
)(
    output reg [COE_WIDTH-1:0] coe0,
    output reg [COE_WIDTH-1:0] coe1,
    output reg [COE_WIDTH-1:0] coe2,
    output reg [COE_WIDTH-1:0] coe3,

    input [$clog2(PIXEL_STEP/4)-1:0] dx,
    input clk
);

(* ROM_STYLE="DISTRIBUTED" *) reg [COE_WIDTH-1:0] coe_table_0[(PIXEL_STEP/4)-1:0];
(* ROM_STYLE="DISTRIBUTED" *) reg [COE_WIDTH-1:0] coe_table_1[(PIXEL_STEP/4)-1:0];
(* ROM_STYLE="DISTRIBUTED" *) reg [COE_WIDTH-1:0] coe_table_2[(PIXEL_STEP/4)-1:0];
(* ROM_STYLE="DISTRIBUTED" *) reg [COE_WIDTH-1:0] coe_table_3[(PIXEL_STEP/4)-1:0];

initial $readmemb("cubic_table_0.txt", coe_table_0);
initial $readmemb("cubic_table_1.txt", coe_table_1);
initial $readmemb("cubic_table_2.txt", coe_table_2);
initial $readmemb("cubic_table_3.txt", coe_table_3);

always @(posedge clk) begin
    coe0 <= coe_table_0[dx];
    coe1 <= coe_table_1[dx];
    coe2 <= coe_table_2[dx];
    coe3 <= coe_table_3[dx];
end

endmodule
