-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 05.06.2012 10:18:05
-- Module Name : video_reader
--
-- ����������/�������� :
--  ������ ����� ����������� �� ���
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_unsigned.all;

library work;
use work.vicg_common_pkg.all;
use work.prj_cfg.all;
use work.prj_def.all;
use work.mem_wr_pkg.all;
use work.dsn_video_ctrl_pkg.all;

entity video_reader is
generic(
G_DBGCS           : string :="OFF";
G_ROTATE          : string:="OFF";
G_ROTATE_BUF_COUNT: integer:=16; --min/max - 4/32
G_MEM_BANK_M_BIT  : integer:=29;
G_MEM_BANK_L_BIT  : integer:=28;

G_MEM_VCH_M_BIT   : integer:=25;
G_MEM_VCH_L_BIT   : integer:=24;
G_MEM_VFR_M_BIT   : integer:=23;
G_MEM_VFR_L_BIT   : integer:=23;
G_MEM_VLINE_M_BIT : integer:=22;
G_MEM_VLINE_L_BIT : integer:=12;

G_MEM_AWIDTH      : integer:=32;
G_MEM_DWIDTH      : integer:=32
);
port(
-------------------------------
-- ����������������
-------------------------------
p_in_cfg_mem_trn_len : in    std_logic_vector(7 downto 0);
p_in_cfg_prm_vch     : in    TReaderVCHParam;

p_in_hrd_chsel       : in    std_logic_vector(3 downto 0);--����: ����� ����������� ��������� ��� ������
p_in_hrd_start       : in    std_logic;                   --����: ������ ������ �����
p_in_hrd_done        : in    std_logic;                   --����: ������������� ������� �����

p_in_vfr_buf         : in    std_logic_vector(G_MEM_VFR_M_BIT - G_MEM_VFR_L_BIT downto 0);
p_in_vfr_nrow        : in    std_logic;                   --���������� ������ ��������� ������

--�������
p_out_vch_fr_new     : out   std_logic;
p_out_vch_rd_done    : out   std_logic;
p_out_vch            : out   std_logic_vector(3 downto 0);
p_out_vch_active_pix : out   std_logic_vector(15 downto 0);
p_out_vch_active_row : out   std_logic_vector(15 downto 0);
p_out_vch_mirx       : out   std_logic;

----------------------------
--Upstream Port
----------------------------
p_out_upp_data       : out   std_logic_vector(G_MEM_DWIDTH - 1 downto 0);
p_out_upp_data_wd    : out   std_logic;
p_in_upp_buf_empty   : in    std_logic;
p_in_upp_buf_full    : in    std_logic;

---------------------------------
-- ����� � mem_ctrl.vhd
---------------------------------
p_out_mem            : out   TMemIN;
p_in_mem             : in    TMemOUT;

-------------------------------
--���������������
-------------------------------
p_in_tst             : in    std_logic_vector(31 downto 0);
p_out_tst            : out   std_logic_vector(31 downto 0);

-------------------------------
--System
-------------------------------
p_in_clk             : in    std_logic;
p_in_rst             : in    std_logic
);
end video_reader;

architecture behavioral of video_reader is

-- Small delay for simulation purposes.
constant dly : time := 1 ps;

type fsm_state is (
S_IDLE,
S_ROW_FINED0,
S_ROW_FINED1,
S_MEM_SET_ADR,
S_MEM_START,
S_MEM_RD,
S_ROW_NXT
);
signal fsm_state_cs: fsm_state;

signal i_mem_ptr                     : std_logic_vector(31 downto 0);
signal i_mem_rdbase                  : std_logic_vector(31 downto 0);
signal i_mem_adr                     : std_logic_vector(31 downto 0);
signal i_mem_trn_len                 : std_logic_vector(15 downto 0);
signal i_mem_dlen_rq                 : std_logic_vector(15 downto 0);
signal i_mem_start                   : std_logic;
signal i_mem_dir                     : std_logic;
signal i_mem_done                    : std_logic;

signal i_vch_num                     : std_logic_vector(p_in_hrd_chsel'high downto 0);
signal i_vfr_mirror                  : TFrXYMirror;
signal i_vfr_row_cnt                 : std_logic_vector(G_MEM_VFR_L_BIT-G_MEM_VLINE_L_BIT downto 0);
signal i_vfr_skip_row                : std_logic_vector(i_vfr_row_cnt'range);
signal i_vfr_active_row              : std_logic_vector(i_vfr_row_cnt'range);
signal i_vfr_done                    : std_logic;
signal i_vfr_new                     : std_logic;
signal i_vfr_buf                     : std_logic_vector(C_VCTRL_MEM_VFR_M_BIT-C_VCTRL_MEM_VFR_L_BIT downto 0);
signal i_vfr_skip_pix                : std_logic_vector(i_vfr_row_cnt'range);
signal i_skip_pix_byte               : std_logic_vector(G_MEM_VLINE_L_BIT - 1 downto 0);
signal i_pix_count_byte              : std_logic_vector(15 downto 0);

signal i_gnd                         : std_logic_vector(G_MEM_DWIDTH - 1 downto 0);

signal tst_fsmstate                  : std_logic_vector(3 downto 0);
signal tst_fsmstate_out              : std_logic_vector(3 downto 0);


--MAIN
begin


------------------------------------
--��������������� �������
------------------------------------
gen_dbgcs_off : if strcmp(G_DBGCS,"OFF") generate
p_out_tst(31 downto 0) <= (others=>'0');
end generate gen_dbgcs_off;

gen_dbgcs_on : if strcmp(G_DBGCS,"ON") generate
p_out_tst(3  downto 0) <= tst_fsmstate_out;
p_out_tst(4)           <= i_mem_start;
p_out_tst(31 downto 5) <= (others=>'0');

process(p_in_clk)
begin
  if rising_edge(p_in_clk) then
    tst_fsmstate_out <= tst_fsmstate;
  end if;
end process;

tst_fsmstate <= CONV_STD_LOGIC_VECTOR(16#02#, tst_fsmstate'length) when fsm_state_cs = S_ROW_FINED0    else
                CONV_STD_LOGIC_VECTOR(16#03#, tst_fsmstate'length) when fsm_state_cs = S_ROW_FINED1    else
                CONV_STD_LOGIC_VECTOR(16#04#, tst_fsmstate'length) when fsm_state_cs = S_MEM_SET_ADR   else
                CONV_STD_LOGIC_VECTOR(16#05#, tst_fsmstate'length) when fsm_state_cs = S_MEM_START     else
                CONV_STD_LOGIC_VECTOR(16#06#, tst_fsmstate'length) when fsm_state_cs = S_MEM_RD        else
                CONV_STD_LOGIC_VECTOR(16#07#, tst_fsmstate'length) when fsm_state_cs = S_ROW_NXT       else
                CONV_STD_LOGIC_VECTOR(16#00#, tst_fsmstate'length); --fsm_state_cs = S_IDLE else
end generate gen_dbgcs_on;

i_gnd <= (others=>'0');


------------------------------------------------
--�������
------------------------------------------------
p_out_vch_rd_done <= i_vfr_done;
p_out_vch_fr_new <= i_vfr_new;

--��������� ������ �������� �����
p_out_vch <= i_vch_num;

p_out_vch_active_pix <= i_pix_count_byte;
p_out_vch_active_row <= EXT(i_vfr_active_row, p_out_vch_active_row'length);
p_out_vch_mirx       <= i_vfr_mirror.pix;


i_vch_num <= p_in_hrd_chsel;

------------------------------------------------
--������� ������ ����� �����
------------------------------------------------
i_pix_count_byte <= p_in_cfg_prm_vch.fr_size.activ.pix(p_in_cfg_prm_vch.fr_size.activ.pix'high - 2 downto 0) & "00";
i_skip_pix_byte <= i_vfr_skip_pix(G_MEM_VLINE_L_BIT - 1 - 2 downto 0) & "00";

--������ ������ ��������
process(p_in_rst,p_in_clk)
  variable vfr_active_row_end : std_logic_vector(i_vfr_row_cnt'range);
begin
  if p_in_rst = '1' then

    fsm_state_cs <= S_IDLE;

    i_mem_rdbase <= (others=>'0');
    i_mem_ptr <= (others=>'0');
    i_mem_adr <= (others=>'0');
    i_mem_trn_len <= (others=>'0');
    i_mem_dlen_rq <= (others=>'0');
    i_mem_dir <= '0';
    i_mem_start <= '0';

    i_vfr_buf <= (others=>'0');
    i_vfr_mirror.pix <= '0';
    i_vfr_mirror.row <= '0';
    i_vfr_row_cnt <= (others=>'0');
    i_vfr_active_row <= (others=>'0');
      vfr_active_row_end := (others=>'0');
    i_vfr_skip_row <= (others=>'0');
    i_vfr_skip_pix <= (others=>'0');

    i_vfr_done <= '0';
    i_vfr_new <= '0';

  elsif rising_edge(p_in_clk) then

    case fsm_state_cs is

      --------------------------------------
      --�������� ���������
      --------------------------------------
      when S_IDLE =>

        i_vfr_done <= '0';

        --�������� ��������� ����� ������
        if p_in_hrd_start = '1' then
          i_mem_trn_len <= EXT(p_in_cfg_mem_trn_len, i_mem_trn_len'length);

          ----------------------------
          --
          ----------------------------
          i_vfr_buf <= p_in_vfr_buf;

          ----------------------------
          --���� ���:
          ----------------------------
          i_mem_rdbase <= p_in_cfg_prm_vch.mem_adr;

          ----------------------------
          --��������������:
          ----------------------------
          i_vfr_mirror.pix <= p_in_cfg_prm_vch.fr_mirror.pix;
          i_vfr_mirror.row <= p_in_cfg_prm_vch.fr_mirror.row;

          ----------------------------
          --�������:
          ----------------------------
          --�������������� ������ ���������� ������
          --(������ ���� ����� ������� ����� ������)
          i_mem_dlen_rq <= EXT(i_pix_count_byte(i_pix_count_byte'high downto log2(G_MEM_DWIDTH/8)), i_mem_dlen_rq'length)
                           + OR_reduce(i_pix_count_byte(log2(G_MEM_DWIDTH/8) - 1 downto 0));

          i_vfr_skip_pix <= p_in_cfg_prm_vch.fr_size.skip.pix(i_vfr_skip_pix'high downto 0);

          ----------------------------
          --������:
          ----------------------------
          i_vfr_active_row <= p_in_cfg_prm_vch.fr_size.activ.row(i_vfr_active_row'high downto 0);
          i_vfr_skip_row <= p_in_cfg_prm_vch.fr_size.skip.row(i_vfr_skip_row'high downto 0);

          --�������������� ������� �����
          if p_in_cfg_prm_vch.fr_mirror.row = '0' then
            i_vfr_row_cnt <= p_in_cfg_prm_vch.fr_size.skip.row(i_vfr_row_cnt'high downto 0);
          else
            i_vfr_row_cnt <= p_in_cfg_prm_vch.fr_size.skip.row(i_vfr_row_cnt'high downto 0)
                             + p_in_cfg_prm_vch.fr_size.activ.row(i_vfr_row_cnt'high downto 0);
          end if;

          i_mem_ptr <= (others=>'0');
          i_vfr_new <= '1';

          fsm_state_cs <= S_ROW_FINED0;
        end if;

      --------------------------------------
      --
      --------------------------------------
      when S_ROW_FINED0 =>

        i_vfr_new <= '0';

        if i_vfr_mirror.row = '1' then
          --�������������� �� Y - ���������
          --�������������� ������� �����
          i_vfr_row_cnt <= i_vfr_row_cnt-1;
        end if;

        vfr_active_row_end := i_vfr_active_row - 1;

        fsm_state_cs <= S_ROW_FINED1;

      --------------------------------------
      --���� ������ ����� �����
      --------------------------------------
      when S_ROW_FINED1 =>

        fsm_state_cs <= S_MEM_SET_ADR;

      --------------------------------------
      --��������� �������� ������ ���
      --------------------------------------
      when S_MEM_SET_ADR =>

        i_mem_ptr(i_mem_ptr'high downto G_MEM_VCH_M_BIT + 1) <= (others=>'0');
        i_mem_ptr(G_MEM_VCH_M_BIT downto G_MEM_VCH_L_BIT) <= i_vch_num(G_MEM_VCH_M_BIT - G_MEM_VCH_L_BIT downto 0);
        i_mem_ptr(G_MEM_VFR_M_BIT downto G_MEM_VFR_L_BIT) <= i_vfr_buf;
        i_mem_ptr(G_MEM_VLINE_M_BIT downto G_MEM_VLINE_L_BIT) <= i_vfr_row_cnt(G_MEM_VLINE_M_BIT - G_MEM_VLINE_L_BIT downto 0);
        i_mem_ptr(G_MEM_VLINE_L_BIT - 1 downto 0) <= i_skip_pix_byte;

        fsm_state_cs <= S_MEM_START;

      --------------------------------------
      --��������� �������� ������ ���
      --------------------------------------
      when S_MEM_START =>

        i_mem_adr <= i_mem_rdbase + i_mem_ptr;
        i_mem_dir <= C_MEMWR_READ;
        i_mem_start <= '1';
        fsm_state_cs <= S_MEM_RD;

      ------------------------------------------------
      --������ ������
      ------------------------------------------------
      when S_MEM_RD =>

        i_mem_start<='0';

        if i_mem_done='1' then
        --�������� ���������
          fsm_state_cs <= S_ROW_NXT;
        end if;

      ------------------------------------------------
      --���� ������� �� ������ ��������� ������
      ------------------------------------------------
      when S_ROW_NXT =>

        if p_in_vfr_nrow = '1' then

          if (i_vfr_mirror.row = '0' and i_vfr_row_cnt = (i_vfr_skip_row + vfr_active_row_end)) or
             (i_vfr_mirror.row = '1' and i_vfr_row_cnt = i_vfr_skip_row) then

              i_vfr_done <= '1';
              fsm_state_cs <= S_IDLE;

          else

            if i_vfr_mirror.row = '1' then
              i_vfr_row_cnt <= i_vfr_row_cnt - 1;
            else
              i_vfr_row_cnt <= i_vfr_row_cnt + 1;
            end if;

            fsm_state_cs <= S_ROW_FINED1;
          end if;

        end if;

    end case;
  end if;
end process;


--------------------------------------------------------
--������ ������/������ ������ ��� (mem_ctrl.vhd)
--------------------------------------------------------
m_mem_wr : mem_wr
generic map(
G_MEM_BANK_M_BIT => G_MEM_BANK_M_BIT,
G_MEM_BANK_L_BIT => G_MEM_BANK_L_BIT,
G_MEM_AWIDTH     => G_MEM_AWIDTH,
G_MEM_DWIDTH     => G_MEM_DWIDTH
)
port map
(
-------------------------------
-- ����������������
-------------------------------
p_in_cfg_mem_adr     => i_mem_adr,
p_in_cfg_mem_trn_len => i_mem_trn_len,
p_in_cfg_mem_dlen_rq => i_mem_dlen_rq,
p_in_cfg_mem_wr      => i_mem_dir,
p_in_cfg_mem_start   => i_mem_start,
p_out_cfg_mem_done   => i_mem_done,

-------------------------------
-- ����� � ����������������� ��������
-------------------------------
p_in_usr_txbuf_dout  => i_gnd,
p_out_usr_txbuf_rd   => open,
p_in_usr_txbuf_empty => '0',

p_out_usr_rxbuf_din  => p_out_upp_data,
p_out_usr_rxbuf_wd   => p_out_upp_data_wd,
p_in_usr_rxbuf_full  => p_in_upp_buf_full,

---------------------------------
-- ����� � mem_ctrl.vhd
---------------------------------
p_out_mem            => p_out_mem,
p_in_mem             => p_in_mem,

-------------------------------
--System
-------------------------------
p_in_tst             => p_in_tst,
p_out_tst            => open,

p_in_clk             => p_in_clk,
p_in_rst             => p_in_rst
);



--END MAIN
end behavioral;


