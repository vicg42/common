-------------------------------------------------------------------------
-- Company     : Linkos
-- Engineer    : Golovachenko Victor
--
-- Create Date : 2010.06
-- Module Name : video_writer
--
-- ����������/�������� :
--  ������ ����� ������������ � ����������� ���
--  � ���������� � ������ �������� ��� ����������� ����� ���
--  ���������������� ����� ������
--
--
-- Revision:
-- Revision 0.01 - File Created
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_unsigned.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.vicg_common_pkg.all;
use work.prj_cfg.all;
use work.prj_def.all;
use work.dsn_video_ctrl_pkg.all;
use work.mem_wr_pkg.all;

entity video_writer is
generic(
G_DBGCS           : string :="OFF";
G_MEM_BANK_M_BIT  : integer:=29;
G_MEM_BANK_L_BIT  : integer:=28;

G_MEM_VCH_M_BIT   : integer:=25;
G_MEM_VCH_L_BIT   : integer:=24;
G_MEM_VFR_M_BIT   : integer:=23;
G_MEM_VFR_L_BIT   : integer:=23;
G_MEM_VLINE_M_BIT : integer:=22;
G_MEM_VLINE_L_BIT : integer:=12;

G_MEM_AWIDTH      : integer:=32;
G_MEM_DWIDTH      : integer:=32
);
port(
-------------------------------
-- ����������������
-------------------------------
p_in_cfg_load         : in    std_logic;                   --//�������� ���������� ������
p_in_cfg_mem_trn_len  : in    std_logic_vector(7 downto 0);--//������ ��������� ���������� MEM_WR
p_in_cfg_prm_vch      : in    TWriterVCHParams;            --//��������� ������ ����� �������
p_in_cfg_set_idle_vch : in    std_logic_vector(C_VCTRL_VCH_COUNT-1 downto 0);

p_in_vfr_buf          : in    TVfrBufs;                    --//����� ������ ��� ����� ������������� ������� ����

--//�������
p_out_vfr_rdy         : out   std_logic_vector(C_VCTRL_VCH_COUNT-1 downto 0);--//���� ����� ��� ���������������� �����������
p_out_vrow_mrk        : out   TVMrks;                      --//������ ������

--//--------------------------
--//Upstream Port (����� � ������� ������������)
--//--------------------------
p_in_upp_data         : in    std_logic_vector(31 downto 0);
p_out_upp_data_rd     : out   std_logic;
p_in_upp_data_rdy     : in    std_logic;
p_in_upp_buf_empty    : in    std_logic;
p_in_upp_buf_full     : in    std_logic;
p_in_upp_buf_pfull    : in    std_logic;

---------------------------------
-- ����� � mem_ctrl.vhd
---------------------------------
p_out_mem             : out   TMemIN;
p_in_mem              : in    TMemOUT;

-------------------------------
--���������������
-------------------------------
p_in_tst              : in    std_logic_vector(31 downto 0);
p_out_tst             : out   std_logic_vector(31 downto 0);

-------------------------------
--System
-------------------------------
p_in_clk              : in    std_logic;
p_in_rst              : in    std_logic
);
end video_writer;

architecture behavioral of video_writer is

-- Small delay for simulation purposes.
constant dly : time := 1 ps;

type fsm_state is (
S_IDLE,
S_PKT_HEADER_READ,
S_MEM_START,
S_MEM_WR,
S_PKT_SKIP
);
signal fsm_state_cs: fsm_state;

signal i_vpkt_cnt                  : std_logic_vector(3 downto 0);
signal i_vpkt_header_rd            : std_logic;
signal i_vpkt_payload_rd           : std_logic;

signal i_vfr_row_mrk               : TVMrks;
signal i_vfr_row_mrk_l             : std_logic_vector(15 downto 0);
signal i_vfr_pix_count             : std_logic_vector(15 downto 0);
signal i_vfr_row_count             : std_logic_vector(15 downto 0);
Type TVfrNum is array (0 to C_VCTRL_VCH_COUNT-1) of std_logic_vector(3 downto 0);
signal i_vfr_num                   : TVfrNum;
signal i_vfr_row                   : std_logic_vector(15 downto 0);
signal i_vch_num                   : std_logic_vector(3 downto 0);
signal i_vfr_rdy                   : std_logic_vector(p_out_vfr_rdy'range);

signal i_mem_ptr                   : std_logic_vector(31 downto 0);
signal i_mem_wrbase                : std_logic_vector(31 downto 0);
signal i_mem_adr                   : std_logic_vector(31 downto 0);
signal i_mem_trn_len               : std_logic_vector(15 downto 0);
signal i_mem_dlen_rq               : std_logic_vector(15 downto 0);
signal i_mem_start                 : std_logic;
signal i_mem_dir                   : std_logic;
signal i_mem_done                  : std_logic;

signal i_upp_data_rd               : std_logic;
signal i_upp_buf_pfull             : std_logic;
signal i_upp_hd_data_rd_out        : std_logic;

signal i_upp_pkt_skip_rd_out       : std_logic;
signal i_pkt_type_err              : std_logic_vector(4 downto 0);
signal i_pkt_size_byte             : std_logic_vector(15 downto 0);
signal i_pkt_size_dw               : std_logic_vector(15 downto 0);
signal i_pkt_sizetotal_byte        : std_logic_vector(15+1 downto 0);
signal i_pkt_skip_dw_calc          : std_logic_vector(15+1+2 downto 0);
signal i_pkt_skip_dw_calc_int      : std_logic_vector(15+1 downto 0);
signal i_pkt_skip_dw_calc_rem      : std_logic_vector(1 downto 0);
signal i_pkt_skip_dw               : std_logic_vector(15+1+1 downto 0);
signal i_pkt_skip_dw_dcnt          : std_logic_vector(15+1+1 downto 0);
signal i_vpkt_size_dw              : std_logic_vector(15 downto 0);
signal i_vpkt_skip_rd              : std_logic;
signal i_vfr_pix_count_dw          : std_logic_vector(15 downto 0);

--signal tst_dbg_pictire             : std_logic;
signal tst_fsmstate                  : std_logic_vector(3 downto 0);
signal tst_fsmstate_out              : std_logic_vector(3 downto 0);
signal tst_upp_buf_empty             : std_logic;


--MAIN
begin


--//----------------------------------
--//��������������� �������
--//----------------------------------
gen_dbgcs_off : if strcmp(G_DBGCS,"OFF") generate
p_out_tst(26 downto 0)<=(others=>'0');
p_out_tst(31 downto 27)<=i_pkt_type_err;
end generate gen_dbgcs_off;

gen_dbgcs_on : if strcmp(G_DBGCS,"ON") generate
p_out_tst(3  downto 0)<=tst_fsmstate_out;
p_out_tst(4)          <=i_mem_start or OR_reduce(i_pkt_type_err) or tst_upp_buf_empty;
p_out_tst(26 downto 5) <=(others=>'0');
p_out_tst(31 downto 27)<=i_pkt_type_err;

process(p_in_clk)
begin
  if p_in_clk'event and p_in_clk='1' then
    tst_fsmstate_out<=tst_fsmstate;
    tst_upp_buf_empty<=p_in_upp_buf_empty;
  end if;
end process;

tst_fsmstate<=CONV_STD_LOGIC_VECTOR(16#01#,tst_fsmstate'length) when fsm_state_cs=S_PKT_HEADER_READ else
              CONV_STD_LOGIC_VECTOR(16#02#,tst_fsmstate'length) when fsm_state_cs=S_MEM_START       else
              CONV_STD_LOGIC_VECTOR(16#03#,tst_fsmstate'length) when fsm_state_cs=S_MEM_WR          else
              CONV_STD_LOGIC_VECTOR(16#04#,tst_fsmstate'length) when fsm_state_cs=S_PKT_SKIP        else
              CONV_STD_LOGIC_VECTOR(16#00#,tst_fsmstate'length); --//fsm_state_cs=S_IDLE              else
end generate gen_dbgcs_on;

--tst_dbg_pictire<=p_in_tst(C_VCTRL_REG_TST0_DBG_PICTURE_BIT);


--//----------------------------------------------
--//�������
--//----------------------------------------------
p_out_vfr_rdy<=i_vfr_rdy;--//����������: ���� ������� � ���
p_out_vrow_mrk<=i_vfr_row_mrk;--//������ ������ ����������


--//----------------------------------------------
--//����� � ������� ����� �������
--//������� ������ ����� ����������
--//----------------------------------------------
p_out_upp_data_rd<=i_upp_hd_data_rd_out or (i_vpkt_payload_rd and i_upp_data_rd) or i_upp_pkt_skip_rd_out;

i_upp_hd_data_rd_out <=(i_vpkt_header_rd  and not p_in_upp_buf_empty);

i_upp_pkt_skip_rd_out <=(i_vpkt_skip_rd  and not p_in_upp_buf_empty);


--//----------------------------------------------
--//
--//----------------------------------------------
--��������� ������� DW ����� ���������� ����� ������� � ������ pkt, ���� �������� ������ � �������� ������
i_pkt_sizetotal_byte<=EXT(i_pkt_size_byte, i_pkt_sizetotal_byte'length) + 2;--���-�� ���� ������ + ���-�� ���� ���� length
i_pkt_skip_dw_calc<="00"&i_pkt_sizetotal_byte(i_pkt_sizetotal_byte'length-1 downto 0);--i_pkt_sizetotal_byte/4
--                                        ����� ����� �� ������� �� 4                              |  ������� �� ������� �� 4
i_pkt_skip_dw<=EXT(i_pkt_skip_dw_calc(i_pkt_skip_dw_calc'length-1 downto 2), i_pkt_skip_dw'length) + OR_reduce(i_pkt_skip_dw_calc(1 downto 0));

--������� ������ ��� ���������
i_vfr_pix_count_dw<=EXT(i_vfr_pix_count(i_vfr_pix_count'high downto 2), i_vfr_pix_count_dw'length) + OR_reduce(i_vfr_pix_count(1 downto 0));
i_vpkt_size_dw<=CONV_STD_LOGIC_VECTOR(C_VIDEO_PKT_HEADER_SIZE, i_vpkt_size_dw'length) + EXT(i_vfr_pix_count_dw, i_vpkt_size_dw'length);
--                                        ����� ����� �� ������� �� 4                        |  ������� �� ������� �� 4
i_pkt_size_dw<=EXT(i_pkt_size_byte(i_pkt_size_byte'length-1 downto 2), i_pkt_size_dw'length) + OR_reduce(i_pkt_size_byte(1 downto 0));

--//----------------------------------------------
--//������� ������ ����� ����������
--//----------------------------------------------
process(p_in_rst,p_in_clk)
  variable vfr_rdy : std_logic_vector(p_out_vfr_rdy'range);
begin
  if p_in_rst='1' then

    fsm_state_cs <= S_IDLE;

    i_vpkt_cnt<=(others=>'0');
    i_vpkt_header_rd<='0';
    i_vpkt_payload_rd<='0';

    i_vch_num<=(others=>'0');
    for i in 0 to C_VCTRL_VCH_COUNT-1 loop
      i_vfr_num(i)<=(others=>'0');
      i_vfr_row_mrk(i)<=(others=>'0');
    end loop;

    i_vfr_row<=(others=>'0');
    i_vfr_pix_count<=(others=>'0');
    i_vfr_row_count<=(others=>'0');
    i_vfr_row_mrk_l<=(others=>'0');
    i_vfr_rdy<=(others=>'0');

    i_upp_buf_pfull<='0';

    vfr_rdy:=(others=>'0');

    i_mem_ptr<=(others=>'0');
    i_mem_wrbase<=(others=>'0');
    i_mem_adr<=(others=>'0');
    i_mem_dlen_rq<=(others=>'0');
    i_mem_trn_len<=(others=>'0');
    i_mem_dir<='0';
    i_mem_start<='0';

    i_vpkt_skip_rd<='0';
    i_pkt_size_byte<=(others=>'0');
    i_pkt_skip_dw_dcnt<=(others=>'0'); i_pkt_type_err<=(others=>'0');

  elsif p_in_clk'event and p_in_clk='1' then

    vfr_rdy:=(others=>'0');

    i_upp_buf_pfull<=p_in_upp_buf_pfull;

    case fsm_state_cs is

      --//------------------------------------
      --//�������� ���������
      --//------------------------------------
      when S_IDLE =>

        i_pkt_skip_dw_dcnt<=(others=>'0'); --i_pkt_type_err<=(others=>'0');

        --//�������� ��������� ����� ������
        if p_in_cfg_load='1' then
          for i in 0 to C_VCTRL_VCH_COUNT-1 loop
            i_mem_wrbase<=p_in_cfg_prm_vch(i).mem_adr;
          end loop;
        end if;

        --//���� ����� �������� ������ � ������
        if i_upp_buf_pfull='1' then --//if p_in_upp_buf_pfull='1' then
        --//���� ����� � ������� ������ ��������� ������ ���-�� ������ (0x40 DWORD)

          i_vpkt_header_rd<='1';
          --//��������� � ������� ������ ��������� ������ ����� ������ (� DWORD)
          i_vpkt_cnt<=CONV_STD_LOGIC_VECTOR(C_VIDEO_PKT_HEADER_SIZE-1, i_vpkt_cnt'length);

          i_pkt_type_err(3 downto 0)<=(others=>'0');
          if p_in_upp_buf_full='1' then
             i_pkt_type_err(4)<='1';
          else
            i_pkt_type_err(4)<='0';
          end if;

          fsm_state_cs <= S_PKT_HEADER_READ;
        end if;

      --//------------------------------------
      --//������ � ������ ��������� ������ �����������
      --//------------------------------------
      when S_PKT_HEADER_READ =>

        if i_upp_hd_data_rd_out='1' then

          i_pkt_skip_dw_dcnt<=i_pkt_skip_dw_dcnt + 1;

          if i_vpkt_cnt=(i_vpkt_cnt'range =>'0') then
          --//----------------------------------------
          --//----- �������� ���� ��������� ----------
          --//----------------------------------------

            i_vpkt_header_rd<='0';

            --//��������� ���������� ��� �������� ����� �����������:
            for i in 0 to C_VCTRL_VCH_COUNT-1 loop
              if i_vch_num=i then

                --//��������� ������ ������� ������ ����� :
                i_vfr_row_mrk(i)(31 downto 16)<=p_in_upp_data(15 downto 0);--//(������� �����)
                i_vfr_row_mrk(i)(15 downto 0)<=i_vfr_row_mrk_l;            --//(������� �����)

                --//����� ���:
                i_mem_ptr(G_MEM_VFR_M_BIT downto G_MEM_VFR_L_BIT)<=p_in_vfr_buf(i);
              end if;
            end loop;

            --//����� ���:
            i_mem_ptr(G_MEM_VCH_M_BIT downto G_MEM_VCH_L_BIT)<=i_vch_num(G_MEM_VCH_M_BIT-G_MEM_VCH_L_BIT downto 0);
            i_mem_ptr(G_MEM_VLINE_M_BIT downto G_MEM_VLINE_L_BIT)<=i_vfr_row((G_MEM_VLINE_M_BIT-G_MEM_VLINE_L_BIT)+0 downto 0);
            i_mem_ptr(G_MEM_VLINE_L_BIT-1 downto 0)<=(others=>'0');--//Pix

            if i_pkt_size_dw=i_vpkt_size_dw then
              fsm_state_cs <= S_MEM_START;
            else
            --Pkt Lenth/4 != (C_VIDEO_PKT_HEADER_SIZE + PIXCOUNT/4)
              i_vpkt_skip_rd<='1'; i_pkt_type_err(3)<='1';
              fsm_state_cs <= S_PKT_SKIP;
            end if;

          else
          --//-------------------------
          --//������ ���������:
          --//-------------------------
            --//Header DWORD-0:
            if i_vpkt_cnt=CONV_STD_LOGIC_VECTOR(C_VIDEO_PKT_HEADER_SIZE-1, i_vpkt_cnt'length) then

              i_pkt_size_byte<=p_in_upp_data(15 downto 0);--Length (byte)

              if p_in_upp_data(19 downto 16)="0001" and p_in_upp_data(27 downto 24)="0011" and p_in_upp_data(23 downto 20)<="0011" then
              --//��� ������ - ����� ������ + �������� ������ ��������� ������

                --//��������� ����� �������� ����� ������:
                i_vch_num<=p_in_upp_data(23 downto 20);
              else
                --//�� ��� �����
                i_vpkt_header_rd<='0';
                i_vpkt_skip_rd<='1';

                if p_in_upp_data(19 downto 16)/="0001" then
                  i_pkt_type_err(0)<='1';--pkt_type
                end if;
                if p_in_upp_data(23 downto 20)>"0011" then
                  i_pkt_type_err(1)<='1';--vch
                end if;
                if p_in_upp_data(27 downto 24)/="0011" then
                  i_pkt_type_err(2)<='1';--src video
                end if;

                fsm_state_cs <= S_PKT_SKIP;
              end if;

            --//Header DWORD-1:
            elsif i_vpkt_cnt=CONV_STD_LOGIC_VECTOR(C_VIDEO_PKT_HEADER_SIZE-2, i_vpkt_cnt'length) then

              for i in 0 to C_VCTRL_VCH_COUNT-1 loop
                if i_vch_num=i then
                  if i_vfr_num(i)/=p_in_upp_data(3 downto 0) then
                    --//��������� ������ ������ �����!!!!!!!!!
                    --//������������ ���������� ������
                    i_mem_wrbase<=p_in_cfg_prm_vch(i).mem_adr;
                  end if;

                  --//��������� ����� �������� �����:
                  i_vfr_num(i)<= p_in_upp_data(3 downto 0);

                 end if;
              end loop;

              --//��������� ������ �����: ���-�� ��������
              i_vfr_pix_count<=p_in_upp_data(31 downto 16);

            --//Header DWORD-2:
            elsif i_vpkt_cnt=CONV_STD_LOGIC_VECTOR(C_VIDEO_PKT_HEADER_SIZE-3, i_vpkt_cnt'length) then

              --//��������� ������ �����: ���-�� �����
              i_vfr_row_count <= p_in_upp_data(15 downto 0);

              --//��������� ����� ������� ������:
              i_vfr_row <= p_in_upp_data(31 downto 16);

            --//Header DWORD-3:
            elsif i_vpkt_cnt=CONV_STD_LOGIC_VECTOR(C_VIDEO_PKT_HEADER_SIZE-4, i_vpkt_cnt'length) then

              --//��������� ������ ������ (������� �����)
              i_vfr_row_mrk_l(15 downto 0)<=p_in_upp_data(31 downto 16);

            end if;

            i_vpkt_cnt<=i_vpkt_cnt-1;

          end if;

        end if;


      --//------------------------------------
      --//��������� �������� ������ ���
      --//------------------------------------
      when S_MEM_START =>

        i_vpkt_payload_rd<='1';
        i_mem_dlen_rq<="00"&i_vfr_pix_count(i_vfr_pix_count'high downto 2); --//DW
        i_mem_trn_len<=EXT(p_in_cfg_mem_trn_len, i_mem_trn_len'length);
        i_mem_adr<=i_mem_wrbase + i_mem_ptr;
        i_mem_dir<=C_MEMWR_WRITE;
        i_mem_start<='1';
        fsm_state_cs <= S_MEM_WR;

      --//----------------------------------------------
      --//������ ������
      --//----------------------------------------------
      when S_MEM_WR =>

        i_mem_start<='0';

        if i_mem_done='1' then
        --//�������� ���������
          i_vpkt_payload_rd<='0';

          if i_vfr_row=(i_vfr_row_count - 1) then
          --//��������� ��������� ������ �����.
          --//������ ����������:
            for i in 0 to C_VCTRL_VCH_COUNT-1 loop
              if i_vch_num=i then
                vfr_rdy(i):='1';
              end if;
            end loop;
          end if;

          fsm_state_cs <= S_IDLE;
        end if;


      --//------------------------------------
      --//������� �������� ������
      --//------------------------------------
      when S_PKT_SKIP =>

        if i_upp_pkt_skip_rd_out='1' then
          if i_pkt_skip_dw_dcnt=(i_pkt_skip_dw - 1) then
            i_vpkt_skip_rd<='0';
            fsm_state_cs <= S_IDLE;
          else
            i_pkt_skip_dw_dcnt<=i_pkt_skip_dw_dcnt + 1;
          end if;
        end if;

    end case;

    i_vfr_rdy<=vfr_rdy;
  end if;
end process;


m_mem_wr : mem_wr
generic map(
G_MEM_BANK_M_BIT => G_MEM_BANK_M_BIT,
G_MEM_BANK_L_BIT => G_MEM_BANK_L_BIT,
G_MEM_AWIDTH     => G_MEM_AWIDTH,
G_MEM_DWIDTH     => G_MEM_DWIDTH
)
port map(
-------------------------------
-- ����������������
-------------------------------
p_in_cfg_mem_adr     => i_mem_adr,
p_in_cfg_mem_trn_len => i_mem_trn_len,
p_in_cfg_mem_dlen_rq => i_mem_dlen_rq,
p_in_cfg_mem_wr      => i_mem_dir,
p_in_cfg_mem_start   => i_mem_start,
p_out_cfg_mem_done   => i_mem_done,

-------------------------------
-- ����� � ����������������� ��������
-------------------------------
p_in_usr_txbuf_dout  => p_in_upp_data,
p_out_usr_txbuf_rd   => i_upp_data_rd,
p_in_usr_txbuf_empty => p_in_upp_buf_empty,

p_out_usr_rxbuf_din  => open,
p_out_usr_rxbuf_wd   => open,
p_in_usr_rxbuf_full  => '0',

---------------------------------
-- ����� � mem_ctrl.vhd
---------------------------------
p_out_mem            => p_out_mem,
p_in_mem             => p_in_mem,

-------------------------------
--System
-------------------------------
p_in_tst             => p_in_tst,
p_out_tst            => open,--tst_mem_ctrl_ch_wr_out,

p_in_clk             => p_in_clk,
p_in_rst             => p_in_rst
);

--END MAIN
end behavioral;

