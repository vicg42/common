//-------------------------------------------------------------
//  ������ ������ � ������� (��������� �����)
//-------------------------------------------------------------
// ����� ������� �.�.
//
// V1.0   6.7.5
// V2.0   31.8.5
// V3.0   22.9.6
//-------------------------------------------------------------
module pult_io(
   input clk_io_en,tmr_en,tmr_stb,             //add vicg
   input rst,clk_io,            //����� � �������� ��� ������ � �������
   input trans_ack,             //���������� PCI �������� ����� � ���-��

   input data_i,                //���������������� ������ �� ������
   output data_o,               //���������������� ������ �� �����
   output dir_485,              //���������� 485 ������-������������

   input host_clk_wr,           //�������� �� ����� ��� ������
   input wr_en,                 //���������� ������ � ������ �����������
   input [31:0] data_from_host, //������ �� ����� ��� ������

   input host_clk_rd,           //�������� �� ����� ��� ������
   input rd_en,                 //���������� ������ � ������ �����������
   output [31:0] data_to_host,  //������ � ����

   output busy,ready           //��������� ������ � �������

);

assign data_o = 0;
assign dir_485 = 0;
assign data_to_host = 0;

assign busy = 0;
assign ready = 0;

endmodule
