//------------------------------------------------------------
// ������ ������������� ����� ������� ���������� ������� ���
//  ������� �����, �������������� ��� ������� ����������������
//  �������� (���� ���������� 3.3���). ����������� ��������
//  ��� �������� �������� ���������������� � ������������� �
//  ���������� �������� �������� �������
// ������ �������: [31]-overday, [30:26]-����, [25:20]-������,
//  [19:14]-�������, [13:4]-��, [3:0]-����� ���.
//------------------------------------------------------------
// ����� ������� �.�.
//
// V1.0     Date 20.4.5 - 24.4.5
// V1.1     Date 14.5.5 - 15.5.5
// V2.0     Date 23.9.6 - 25.9.6
// V2.1     Date 24.10.6 - 24.10.6
// V2.2     Date 2.11.6
// V2.3     Date 30.06.10 ������� ���� ������� ��� ������������������� ���������
//------------------------- -----------------------------------
module sync_u(
   input i_clk,
   input i_pps,i_ext_1s,i_ext_1m,		 //PPS � ������� �������������

   input sync_iedge,       //����������� ������ ������ ������� ������������� (0-rise)
   input sync_oedge,       //����������� ������ ������� �� ������� ������������� (0-rise)
   input sync_time_en,     //���������� ������ ����� (1-���������)
   input mode_set_time,    //��������� ����� (0-����� � �������, 1-�� ������� �������)
   input [1:0] type_of_sync, //����� ��������� ������� �������������,
// '10'-�������, '01'-PPS, '11','00'-���������� �������������

   output sync_win,         //���������� �������� ������ ������� (1 ��)

   input host_clk,               //�������� �� �����
   input wr_en_time,             //��������� �������
   input [31:0] host_wr_data,   //������ �� ����� ��� ������

   output [31:0] stime,          //���������� ������� �������
   output [7:0] n_sync,          //����� ��������������
   output [7:0] sync_cou_err,    //������� ������ ������� ������������� (�� � �������)

   output sync_out1,out_1s,out_1m,    //������������� ��� ������� ���������
	output sync_out2,
	output sync_ld,  //������������� ��
	output sync_pic  //������������� PIC
);


assign sync_win = 0;

assign stime = 0;
assign n_sync = 0;
assign sync_cou_err = 0;

assign sync_out1 = 0;
assign out_1s = 0;
assign out_1m = 0;
assign sync_out2 = 0;
assign sync_ld = 0;
assign sync_pic = 0;

endmodule
